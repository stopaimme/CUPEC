`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/09/25 15:31:14
// Design Name: 
// Module Name: ultra
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ultra(
    input clk,
    input reset,
    output reg [24:0] io0,
output reg [24:0] io1,
output reg [24:0] io2,
output reg [24:0] io3,
output reg [24:0] io4,
output reg [24:0] io5,
output reg [24:0] io6,
output reg [24:0] io7,
output reg [24:0] io8,
output reg [24:0] io9,
output reg [24:0] io10,
output reg [24:0] io11,
output reg [24:0] io12,
output reg [24:0] io13,
output reg [24:0] io14,
output reg [24:0] io15,
output reg [24:0] io16,
output reg [24:0] io17,
output reg [24:0] io18,
output reg [24:0] io19,
output reg [24:0] io20,
output reg [24:0] io21,
output reg [24:0] io22,
output reg [24:0] io23,
output reg [24:0] io24,
output reg [24:0] io25,
output reg [24:0] io26,
output reg [24:0] io27,
output reg [24:0] io28,
output reg [24:0] io29,
output reg [24:0] io30,
output reg [24:0] io31,
output reg [24:0] io32,
output reg [24:0] io33,
output reg [24:0] io34,
output reg [24:0] io35,
output reg [24:0] io36,
output reg [24:0] io37,
output reg [24:0] io38,
output reg [24:0] io39
    );
reg [10:0] m0_0;
reg [10:0] m0_1;
reg [10:0] m0_2;
reg [10:0] m0_3;
reg [10:0] m0_4;
reg [10:0] m0_5;
reg [10:0] m0_6;
reg [10:0] m0_7;
reg [10:0] m0_8;
reg [10:0] m0_9;
reg [10:0] m0_10;
reg [10:0] m0_11;
reg [10:0] m0_12;
reg [10:0] m0_13;
reg [10:0] m0_14;
reg [10:0] m0_15;
reg [10:0] m0_16;
reg [10:0] m0_17;
reg [10:0] m0_18;
reg [10:0] m0_19;
reg [10:0] m0_20;
reg [10:0] m0_21;
reg [10:0] m0_22;
reg [10:0] m0_23;
reg [10:0] m0_24;
reg [10:0] m1_0;
reg [10:0] m1_1;
reg [10:0] m1_2;
reg [10:0] m1_3;
reg [10:0] m1_4;
reg [10:0] m1_5;
reg [10:0] m1_6;
reg [10:0] m1_7;
reg [10:0] m1_8;
reg [10:0] m1_9;
reg [10:0] m1_10;
reg [10:0] m1_11;
reg [10:0] m1_12;
reg [10:0] m1_13;
reg [10:0] m1_14;
reg [10:0] m1_15;
reg [10:0] m1_16;
reg [10:0] m1_17;
reg [10:0] m1_18;
reg [10:0] m1_19;
reg [10:0] m1_20;
reg [10:0] m1_21;
reg [10:0] m1_22;
reg [10:0] m1_23;
reg [10:0] m1_24;
reg [10:0] m2_0;
reg [10:0] m2_1;
reg [10:0] m2_2;
reg [10:0] m2_3;
reg [10:0] m2_4;
reg [10:0] m2_5;
reg [10:0] m2_6;
reg [10:0] m2_7;
reg [10:0] m2_8;
reg [10:0] m2_9;
reg [10:0] m2_10;
reg [10:0] m2_11;
reg [10:0] m2_12;
reg [10:0] m2_13;
reg [10:0] m2_14;
reg [10:0] m2_15;
reg [10:0] m2_16;
reg [10:0] m2_17;
reg [10:0] m2_18;
reg [10:0] m2_19;
reg [10:0] m2_20;
reg [10:0] m2_21;
reg [10:0] m2_22;
reg [10:0] m2_23;
reg [10:0] m2_24;
reg [10:0] m3_0;
reg [10:0] m3_1;
reg [10:0] m3_2;
reg [10:0] m3_3;
reg [10:0] m3_4;
reg [10:0] m3_5;
reg [10:0] m3_6;
reg [10:0] m3_7;
reg [10:0] m3_8;
reg [10:0] m3_9;
reg [10:0] m3_10;
reg [10:0] m3_11;
reg [10:0] m3_12;
reg [10:0] m3_13;
reg [10:0] m3_14;
reg [10:0] m3_15;
reg [10:0] m3_16;
reg [10:0] m3_17;
reg [10:0] m3_18;
reg [10:0] m3_19;
reg [10:0] m3_20;
reg [10:0] m3_21;
reg [10:0] m3_22;
reg [10:0] m3_23;
reg [10:0] m3_24;
reg [10:0] m4_0;
reg [10:0] m4_1;
reg [10:0] m4_2;
reg [10:0] m4_3;
reg [10:0] m4_4;
reg [10:0] m4_5;
reg [10:0] m4_6;
reg [10:0] m4_7;
reg [10:0] m4_8;
reg [10:0] m4_9;
reg [10:0] m4_10;
reg [10:0] m4_11;
reg [10:0] m4_12;
reg [10:0] m4_13;
reg [10:0] m4_14;
reg [10:0] m4_15;
reg [10:0] m4_16;
reg [10:0] m4_17;
reg [10:0] m4_18;
reg [10:0] m4_19;
reg [10:0] m4_20;
reg [10:0] m4_21;
reg [10:0] m4_22;
reg [10:0] m4_23;
reg [10:0] m4_24;
reg [10:0] m5_0;
reg [10:0] m5_1;
reg [10:0] m5_2;
reg [10:0] m5_3;
reg [10:0] m5_4;
reg [10:0] m5_5;
reg [10:0] m5_6;
reg [10:0] m5_7;
reg [10:0] m5_8;
reg [10:0] m5_9;
reg [10:0] m5_10;
reg [10:0] m5_11;
reg [10:0] m5_12;
reg [10:0] m5_13;
reg [10:0] m5_14;
reg [10:0] m5_15;
reg [10:0] m5_16;
reg [10:0] m5_17;
reg [10:0] m5_18;
reg [10:0] m5_19;
reg [10:0] m5_20;
reg [10:0] m5_21;
reg [10:0] m5_22;
reg [10:0] m5_23;
reg [10:0] m5_24;
reg [10:0] m6_0;
reg [10:0] m6_1;
reg [10:0] m6_2;
reg [10:0] m6_3;
reg [10:0] m6_4;
reg [10:0] m6_5;
reg [10:0] m6_6;
reg [10:0] m6_7;
reg [10:0] m6_8;
reg [10:0] m6_9;
reg [10:0] m6_10;
reg [10:0] m6_11;
reg [10:0] m6_12;
reg [10:0] m6_13;
reg [10:0] m6_14;
reg [10:0] m6_15;
reg [10:0] m6_16;
reg [10:0] m6_17;
reg [10:0] m6_18;
reg [10:0] m6_19;
reg [10:0] m6_20;
reg [10:0] m6_21;
reg [10:0] m6_22;
reg [10:0] m6_23;
reg [10:0] m6_24;
reg [10:0] m7_0;
reg [10:0] m7_1;
reg [10:0] m7_2;
reg [10:0] m7_3;
reg [10:0] m7_4;
reg [10:0] m7_5;
reg [10:0] m7_6;
reg [10:0] m7_7;
reg [10:0] m7_8;
reg [10:0] m7_9;
reg [10:0] m7_10;
reg [10:0] m7_11;
reg [10:0] m7_12;
reg [10:0] m7_13;
reg [10:0] m7_14;
reg [10:0] m7_15;
reg [10:0] m7_16;
reg [10:0] m7_17;
reg [10:0] m7_18;
reg [10:0] m7_19;
reg [10:0] m7_20;
reg [10:0] m7_21;
reg [10:0] m7_22;
reg [10:0] m7_23;
reg [10:0] m7_24;
reg [10:0] m8_0;
reg [10:0] m8_1;
reg [10:0] m8_2;
reg [10:0] m8_3;
reg [10:0] m8_4;
reg [10:0] m8_5;
reg [10:0] m8_6;
reg [10:0] m8_7;
reg [10:0] m8_8;
reg [10:0] m8_9;
reg [10:0] m8_10;
reg [10:0] m8_11;
reg [10:0] m8_12;
reg [10:0] m8_13;
reg [10:0] m8_14;
reg [10:0] m8_15;
reg [10:0] m8_16;
reg [10:0] m8_17;
reg [10:0] m8_18;
reg [10:0] m8_19;
reg [10:0] m8_20;
reg [10:0] m8_21;
reg [10:0] m8_22;
reg [10:0] m8_23;
reg [10:0] m8_24;
reg [10:0] m9_0;
reg [10:0] m9_1;
reg [10:0] m9_2;
reg [10:0] m9_3;
reg [10:0] m9_4;
reg [10:0] m9_5;
reg [10:0] m9_6;
reg [10:0] m9_7;
reg [10:0] m9_8;
reg [10:0] m9_9;
reg [10:0] m9_10;
reg [10:0] m9_11;
reg [10:0] m9_12;
reg [10:0] m9_13;
reg [10:0] m9_14;
reg [10:0] m9_15;
reg [10:0] m9_16;
reg [10:0] m9_17;
reg [10:0] m9_18;
reg [10:0] m9_19;
reg [10:0] m9_20;
reg [10:0] m9_21;
reg [10:0] m9_22;
reg [10:0] m9_23;
reg [10:0] m9_24;
reg [10:0] m10_0;
reg [10:0] m10_1;
reg [10:0] m10_2;
reg [10:0] m10_3;
reg [10:0] m10_4;
reg [10:0] m10_5;
reg [10:0] m10_6;
reg [10:0] m10_7;
reg [10:0] m10_8;
reg [10:0] m10_9;
reg [10:0] m10_10;
reg [10:0] m10_11;
reg [10:0] m10_12;
reg [10:0] m10_13;
reg [10:0] m10_14;
reg [10:0] m10_15;
reg [10:0] m10_16;
reg [10:0] m10_17;
reg [10:0] m10_18;
reg [10:0] m10_19;
reg [10:0] m10_20;
reg [10:0] m10_21;
reg [10:0] m10_22;
reg [10:0] m10_23;
reg [10:0] m10_24;
reg [10:0] m11_0;
reg [10:0] m11_1;
reg [10:0] m11_2;
reg [10:0] m11_3;
reg [10:0] m11_4;
reg [10:0] m11_5;
reg [10:0] m11_6;
reg [10:0] m11_7;
reg [10:0] m11_8;
reg [10:0] m11_9;
reg [10:0] m11_10;
reg [10:0] m11_11;
reg [10:0] m11_12;
reg [10:0] m11_13;
reg [10:0] m11_14;
reg [10:0] m11_15;
reg [10:0] m11_16;
reg [10:0] m11_17;
reg [10:0] m11_18;
reg [10:0] m11_19;
reg [10:0] m11_20;
reg [10:0] m11_21;
reg [10:0] m11_22;
reg [10:0] m11_23;
reg [10:0] m11_24;
reg [10:0] m12_0;
reg [10:0] m12_1;
reg [10:0] m12_2;
reg [10:0] m12_3;
reg [10:0] m12_4;
reg [10:0] m12_5;
reg [10:0] m12_6;
reg [10:0] m12_7;
reg [10:0] m12_8;
reg [10:0] m12_9;
reg [10:0] m12_10;
reg [10:0] m12_11;
reg [10:0] m12_12;
reg [10:0] m12_13;
reg [10:0] m12_14;
reg [10:0] m12_15;
reg [10:0] m12_16;
reg [10:0] m12_17;
reg [10:0] m12_18;
reg [10:0] m12_19;
reg [10:0] m12_20;
reg [10:0] m12_21;
reg [10:0] m12_22;
reg [10:0] m12_23;
reg [10:0] m12_24;
reg [10:0] m13_0;
reg [10:0] m13_1;
reg [10:0] m13_2;
reg [10:0] m13_3;
reg [10:0] m13_4;
reg [10:0] m13_5;
reg [10:0] m13_6;
reg [10:0] m13_7;
reg [10:0] m13_8;
reg [10:0] m13_9;
reg [10:0] m13_10;
reg [10:0] m13_11;
reg [10:0] m13_12;
reg [10:0] m13_13;
reg [10:0] m13_14;
reg [10:0] m13_15;
reg [10:0] m13_16;
reg [10:0] m13_17;
reg [10:0] m13_18;
reg [10:0] m13_19;
reg [10:0] m13_20;
reg [10:0] m13_21;
reg [10:0] m13_22;
reg [10:0] m13_23;
reg [10:0] m13_24;
reg [10:0] m14_0;
reg [10:0] m14_1;
reg [10:0] m14_2;
reg [10:0] m14_3;
reg [10:0] m14_4;
reg [10:0] m14_5;
reg [10:0] m14_6;
reg [10:0] m14_7;
reg [10:0] m14_8;
reg [10:0] m14_9;
reg [10:0] m14_10;
reg [10:0] m14_11;
reg [10:0] m14_12;
reg [10:0] m14_13;
reg [10:0] m14_14;
reg [10:0] m14_15;
reg [10:0] m14_16;
reg [10:0] m14_17;
reg [10:0] m14_18;
reg [10:0] m14_19;
reg [10:0] m14_20;
reg [10:0] m14_21;
reg [10:0] m14_22;
reg [10:0] m14_23;
reg [10:0] m14_24;
reg [10:0] m15_0;
reg [10:0] m15_1;
reg [10:0] m15_2;
reg [10:0] m15_3;
reg [10:0] m15_4;
reg [10:0] m15_5;
reg [10:0] m15_6;
reg [10:0] m15_7;
reg [10:0] m15_8;
reg [10:0] m15_9;
reg [10:0] m15_10;
reg [10:0] m15_11;
reg [10:0] m15_12;
reg [10:0] m15_13;
reg [10:0] m15_14;
reg [10:0] m15_15;
reg [10:0] m15_16;
reg [10:0] m15_17;
reg [10:0] m15_18;
reg [10:0] m15_19;
reg [10:0] m15_20;
reg [10:0] m15_21;
reg [10:0] m15_22;
reg [10:0] m15_23;
reg [10:0] m15_24;
reg [10:0] m16_0;
reg [10:0] m16_1;
reg [10:0] m16_2;
reg [10:0] m16_3;
reg [10:0] m16_4;
reg [10:0] m16_5;
reg [10:0] m16_6;
reg [10:0] m16_7;
reg [10:0] m16_8;
reg [10:0] m16_9;
reg [10:0] m16_10;
reg [10:0] m16_11;
reg [10:0] m16_12;
reg [10:0] m16_13;
reg [10:0] m16_14;
reg [10:0] m16_15;
reg [10:0] m16_16;
reg [10:0] m16_17;
reg [10:0] m16_18;
reg [10:0] m16_19;
reg [10:0] m16_20;
reg [10:0] m16_21;
reg [10:0] m16_22;
reg [10:0] m16_23;
reg [10:0] m16_24;
reg [10:0] m17_0;
reg [10:0] m17_1;
reg [10:0] m17_2;
reg [10:0] m17_3;
reg [10:0] m17_4;
reg [10:0] m17_5;
reg [10:0] m17_6;
reg [10:0] m17_7;
reg [10:0] m17_8;
reg [10:0] m17_9;
reg [10:0] m17_10;
reg [10:0] m17_11;
reg [10:0] m17_12;
reg [10:0] m17_13;
reg [10:0] m17_14;
reg [10:0] m17_15;
reg [10:0] m17_16;
reg [10:0] m17_17;
reg [10:0] m17_18;
reg [10:0] m17_19;
reg [10:0] m17_20;
reg [10:0] m17_21;
reg [10:0] m17_22;
reg [10:0] m17_23;
reg [10:0] m17_24;
reg [10:0] m18_0;
reg [10:0] m18_1;
reg [10:0] m18_2;
reg [10:0] m18_3;
reg [10:0] m18_4;
reg [10:0] m18_5;
reg [10:0] m18_6;
reg [10:0] m18_7;
reg [10:0] m18_8;
reg [10:0] m18_9;
reg [10:0] m18_10;
reg [10:0] m18_11;
reg [10:0] m18_12;
reg [10:0] m18_13;
reg [10:0] m18_14;
reg [10:0] m18_15;
reg [10:0] m18_16;
reg [10:0] m18_17;
reg [10:0] m18_18;
reg [10:0] m18_19;
reg [10:0] m18_20;
reg [10:0] m18_21;
reg [10:0] m18_22;
reg [10:0] m18_23;
reg [10:0] m18_24;
reg [10:0] m19_0;
reg [10:0] m19_1;
reg [10:0] m19_2;
reg [10:0] m19_3;
reg [10:0] m19_4;
reg [10:0] m19_5;
reg [10:0] m19_6;
reg [10:0] m19_7;
reg [10:0] m19_8;
reg [10:0] m19_9;
reg [10:0] m19_10;
reg [10:0] m19_11;
reg [10:0] m19_12;
reg [10:0] m19_13;
reg [10:0] m19_14;
reg [10:0] m19_15;
reg [10:0] m19_16;
reg [10:0] m19_17;
reg [10:0] m19_18;
reg [10:0] m19_19;
reg [10:0] m19_20;
reg [10:0] m19_21;
reg [10:0] m19_22;
reg [10:0] m19_23;
reg [10:0] m19_24;
reg [10:0] m20_0;
reg [10:0] m20_1;
reg [10:0] m20_2;
reg [10:0] m20_3;
reg [10:0] m20_4;
reg [10:0] m20_5;
reg [10:0] m20_6;
reg [10:0] m20_7;
reg [10:0] m20_8;
reg [10:0] m20_9;
reg [10:0] m20_10;
reg [10:0] m20_11;
reg [10:0] m20_12;
reg [10:0] m20_13;
reg [10:0] m20_14;
reg [10:0] m20_15;
reg [10:0] m20_16;
reg [10:0] m20_17;
reg [10:0] m20_18;
reg [10:0] m20_19;
reg [10:0] m20_20;
reg [10:0] m20_21;
reg [10:0] m20_22;
reg [10:0] m20_23;
reg [10:0] m20_24;
reg [10:0] m21_0;
reg [10:0] m21_1;
reg [10:0] m21_2;
reg [10:0] m21_3;
reg [10:0] m21_4;
reg [10:0] m21_5;
reg [10:0] m21_6;
reg [10:0] m21_7;
reg [10:0] m21_8;
reg [10:0] m21_9;
reg [10:0] m21_10;
reg [10:0] m21_11;
reg [10:0] m21_12;
reg [10:0] m21_13;
reg [10:0] m21_14;
reg [10:0] m21_15;
reg [10:0] m21_16;
reg [10:0] m21_17;
reg [10:0] m21_18;
reg [10:0] m21_19;
reg [10:0] m21_20;
reg [10:0] m21_21;
reg [10:0] m21_22;
reg [10:0] m21_23;
reg [10:0] m21_24;
reg [10:0] m22_0;
reg [10:0] m22_1;
reg [10:0] m22_2;
reg [10:0] m22_3;
reg [10:0] m22_4;
reg [10:0] m22_5;
reg [10:0] m22_6;
reg [10:0] m22_7;
reg [10:0] m22_8;
reg [10:0] m22_9;
reg [10:0] m22_10;
reg [10:0] m22_11;
reg [10:0] m22_12;
reg [10:0] m22_13;
reg [10:0] m22_14;
reg [10:0] m22_15;
reg [10:0] m22_16;
reg [10:0] m22_17;
reg [10:0] m22_18;
reg [10:0] m22_19;
reg [10:0] m22_20;
reg [10:0] m22_21;
reg [10:0] m22_22;
reg [10:0] m22_23;
reg [10:0] m22_24;
reg [10:0] m23_0;
reg [10:0] m23_1;
reg [10:0] m23_2;
reg [10:0] m23_3;
reg [10:0] m23_4;
reg [10:0] m23_5;
reg [10:0] m23_6;
reg [10:0] m23_7;
reg [10:0] m23_8;
reg [10:0] m23_9;
reg [10:0] m23_10;
reg [10:0] m23_11;
reg [10:0] m23_12;
reg [10:0] m23_13;
reg [10:0] m23_14;
reg [10:0] m23_15;
reg [10:0] m23_16;
reg [10:0] m23_17;
reg [10:0] m23_18;
reg [10:0] m23_19;
reg [10:0] m23_20;
reg [10:0] m23_21;
reg [10:0] m23_22;
reg [10:0] m23_23;
reg [10:0] m23_24;
reg [10:0] m24_0;
reg [10:0] m24_1;
reg [10:0] m24_2;
reg [10:0] m24_3;
reg [10:0] m24_4;
reg [10:0] m24_5;
reg [10:0] m24_6;
reg [10:0] m24_7;
reg [10:0] m24_8;
reg [10:0] m24_9;
reg [10:0] m24_10;
reg [10:0] m24_11;
reg [10:0] m24_12;
reg [10:0] m24_13;
reg [10:0] m24_14;
reg [10:0] m24_15;
reg [10:0] m24_16;
reg [10:0] m24_17;
reg [10:0] m24_18;
reg [10:0] m24_19;
reg [10:0] m24_20;
reg [10:0] m24_21;
reg [10:0] m24_22;
reg [10:0] m24_23;
reg [10:0] m24_24;
reg [10:0] m25_0;
reg [10:0] m25_1;
reg [10:0] m25_2;
reg [10:0] m25_3;
reg [10:0] m25_4;
reg [10:0] m25_5;
reg [10:0] m25_6;
reg [10:0] m25_7;
reg [10:0] m25_8;
reg [10:0] m25_9;
reg [10:0] m25_10;
reg [10:0] m25_11;
reg [10:0] m25_12;
reg [10:0] m25_13;
reg [10:0] m25_14;
reg [10:0] m25_15;
reg [10:0] m25_16;
reg [10:0] m25_17;
reg [10:0] m25_18;
reg [10:0] m25_19;
reg [10:0] m25_20;
reg [10:0] m25_21;
reg [10:0] m25_22;
reg [10:0] m25_23;
reg [10:0] m25_24;
reg [10:0] m26_0;
reg [10:0] m26_1;
reg [10:0] m26_2;
reg [10:0] m26_3;
reg [10:0] m26_4;
reg [10:0] m26_5;
reg [10:0] m26_6;
reg [10:0] m26_7;
reg [10:0] m26_8;
reg [10:0] m26_9;
reg [10:0] m26_10;
reg [10:0] m26_11;
reg [10:0] m26_12;
reg [10:0] m26_13;
reg [10:0] m26_14;
reg [10:0] m26_15;
reg [10:0] m26_16;
reg [10:0] m26_17;
reg [10:0] m26_18;
reg [10:0] m26_19;
reg [10:0] m26_20;
reg [10:0] m26_21;
reg [10:0] m26_22;
reg [10:0] m26_23;
reg [10:0] m26_24;
reg [10:0] m27_0;
reg [10:0] m27_1;
reg [10:0] m27_2;
reg [10:0] m27_3;
reg [10:0] m27_4;
reg [10:0] m27_5;
reg [10:0] m27_6;
reg [10:0] m27_7;
reg [10:0] m27_8;
reg [10:0] m27_9;
reg [10:0] m27_10;
reg [10:0] m27_11;
reg [10:0] m27_12;
reg [10:0] m27_13;
reg [10:0] m27_14;
reg [10:0] m27_15;
reg [10:0] m27_16;
reg [10:0] m27_17;
reg [10:0] m27_18;
reg [10:0] m27_19;
reg [10:0] m27_20;
reg [10:0] m27_21;
reg [10:0] m27_22;
reg [10:0] m27_23;
reg [10:0] m27_24;
reg [10:0] m28_0;
reg [10:0] m28_1;
reg [10:0] m28_2;
reg [10:0] m28_3;
reg [10:0] m28_4;
reg [10:0] m28_5;
reg [10:0] m28_6;
reg [10:0] m28_7;
reg [10:0] m28_8;
reg [10:0] m28_9;
reg [10:0] m28_10;
reg [10:0] m28_11;
reg [10:0] m28_12;
reg [10:0] m28_13;
reg [10:0] m28_14;
reg [10:0] m28_15;
reg [10:0] m28_16;
reg [10:0] m28_17;
reg [10:0] m28_18;
reg [10:0] m28_19;
reg [10:0] m28_20;
reg [10:0] m28_21;
reg [10:0] m28_22;
reg [10:0] m28_23;
reg [10:0] m28_24;
reg [10:0] m29_0;
reg [10:0] m29_1;
reg [10:0] m29_2;
reg [10:0] m29_3;
reg [10:0] m29_4;
reg [10:0] m29_5;
reg [10:0] m29_6;
reg [10:0] m29_7;
reg [10:0] m29_8;
reg [10:0] m29_9;
reg [10:0] m29_10;
reg [10:0] m29_11;
reg [10:0] m29_12;
reg [10:0] m29_13;
reg [10:0] m29_14;
reg [10:0] m29_15;
reg [10:0] m29_16;
reg [10:0] m29_17;
reg [10:0] m29_18;
reg [10:0] m29_19;
reg [10:0] m29_20;
reg [10:0] m29_21;
reg [10:0] m29_22;
reg [10:0] m29_23;
reg [10:0] m29_24;
reg [10:0] m30_0;
reg [10:0] m30_1;
reg [10:0] m30_2;
reg [10:0] m30_3;
reg [10:0] m30_4;
reg [10:0] m30_5;
reg [10:0] m30_6;
reg [10:0] m30_7;
reg [10:0] m30_8;
reg [10:0] m30_9;
reg [10:0] m30_10;
reg [10:0] m30_11;
reg [10:0] m30_12;
reg [10:0] m30_13;
reg [10:0] m30_14;
reg [10:0] m30_15;
reg [10:0] m30_16;
reg [10:0] m30_17;
reg [10:0] m30_18;
reg [10:0] m30_19;
reg [10:0] m30_20;
reg [10:0] m30_21;
reg [10:0] m30_22;
reg [10:0] m30_23;
reg [10:0] m30_24;
reg [10:0] m31_0;
reg [10:0] m31_1;
reg [10:0] m31_2;
reg [10:0] m31_3;
reg [10:0] m31_4;
reg [10:0] m31_5;
reg [10:0] m31_6;
reg [10:0] m31_7;
reg [10:0] m31_8;
reg [10:0] m31_9;
reg [10:0] m31_10;
reg [10:0] m31_11;
reg [10:0] m31_12;
reg [10:0] m31_13;
reg [10:0] m31_14;
reg [10:0] m31_15;
reg [10:0] m31_16;
reg [10:0] m31_17;
reg [10:0] m31_18;
reg [10:0] m31_19;
reg [10:0] m31_20;
reg [10:0] m31_21;
reg [10:0] m31_22;
reg [10:0] m31_23;
reg [10:0] m31_24;
reg [10:0] m32_0;
reg [10:0] m32_1;
reg [10:0] m32_2;
reg [10:0] m32_3;
reg [10:0] m32_4;
reg [10:0] m32_5;
reg [10:0] m32_6;
reg [10:0] m32_7;
reg [10:0] m32_8;
reg [10:0] m32_9;
reg [10:0] m32_10;
reg [10:0] m32_11;
reg [10:0] m32_12;
reg [10:0] m32_13;
reg [10:0] m32_14;
reg [10:0] m32_15;
reg [10:0] m32_16;
reg [10:0] m32_17;
reg [10:0] m32_18;
reg [10:0] m32_19;
reg [10:0] m32_20;
reg [10:0] m32_21;
reg [10:0] m32_22;
reg [10:0] m32_23;
reg [10:0] m32_24;
reg [10:0] m33_0;
reg [10:0] m33_1;
reg [10:0] m33_2;
reg [10:0] m33_3;
reg [10:0] m33_4;
reg [10:0] m33_5;
reg [10:0] m33_6;
reg [10:0] m33_7;
reg [10:0] m33_8;
reg [10:0] m33_9;
reg [10:0] m33_10;
reg [10:0] m33_11;
reg [10:0] m33_12;
reg [10:0] m33_13;
reg [10:0] m33_14;
reg [10:0] m33_15;
reg [10:0] m33_16;
reg [10:0] m33_17;
reg [10:0] m33_18;
reg [10:0] m33_19;
reg [10:0] m33_20;
reg [10:0] m33_21;
reg [10:0] m33_22;
reg [10:0] m33_23;
reg [10:0] m33_24;
reg [10:0] m34_0;
reg [10:0] m34_1;
reg [10:0] m34_2;
reg [10:0] m34_3;
reg [10:0] m34_4;
reg [10:0] m34_5;
reg [10:0] m34_6;
reg [10:0] m34_7;
reg [10:0] m34_8;
reg [10:0] m34_9;
reg [10:0] m34_10;
reg [10:0] m34_11;
reg [10:0] m34_12;
reg [10:0] m34_13;
reg [10:0] m34_14;
reg [10:0] m34_15;
reg [10:0] m34_16;
reg [10:0] m34_17;
reg [10:0] m34_18;
reg [10:0] m34_19;
reg [10:0] m34_20;
reg [10:0] m34_21;
reg [10:0] m34_22;
reg [10:0] m34_23;
reg [10:0] m34_24;
reg [10:0] m35_0;
reg [10:0] m35_1;
reg [10:0] m35_2;
reg [10:0] m35_3;
reg [10:0] m35_4;
reg [10:0] m35_5;
reg [10:0] m35_6;
reg [10:0] m35_7;
reg [10:0] m35_8;
reg [10:0] m35_9;
reg [10:0] m35_10;
reg [10:0] m35_11;
reg [10:0] m35_12;
reg [10:0] m35_13;
reg [10:0] m35_14;
reg [10:0] m35_15;
reg [10:0] m35_16;
reg [10:0] m35_17;
reg [10:0] m35_18;
reg [10:0] m35_19;
reg [10:0] m35_20;
reg [10:0] m35_21;
reg [10:0] m35_22;
reg [10:0] m35_23;
reg [10:0] m35_24;
reg [10:0] m36_0;
reg [10:0] m36_1;
reg [10:0] m36_2;
reg [10:0] m36_3;
reg [10:0] m36_4;
reg [10:0] m36_5;
reg [10:0] m36_6;
reg [10:0] m36_7;
reg [10:0] m36_8;
reg [10:0] m36_9;
reg [10:0] m36_10;
reg [10:0] m36_11;
reg [10:0] m36_12;
reg [10:0] m36_13;
reg [10:0] m36_14;
reg [10:0] m36_15;
reg [10:0] m36_16;
reg [10:0] m36_17;
reg [10:0] m36_18;
reg [10:0] m36_19;
reg [10:0] m36_20;
reg [10:0] m36_21;
reg [10:0] m36_22;
reg [10:0] m36_23;
reg [10:0] m36_24;
reg [10:0] m37_0;
reg [10:0] m37_1;
reg [10:0] m37_2;
reg [10:0] m37_3;
reg [10:0] m37_4;
reg [10:0] m37_5;
reg [10:0] m37_6;
reg [10:0] m37_7;
reg [10:0] m37_8;
reg [10:0] m37_9;
reg [10:0] m37_10;
reg [10:0] m37_11;
reg [10:0] m37_12;
reg [10:0] m37_13;
reg [10:0] m37_14;
reg [10:0] m37_15;
reg [10:0] m37_16;
reg [10:0] m37_17;
reg [10:0] m37_18;
reg [10:0] m37_19;
reg [10:0] m37_20;
reg [10:0] m37_21;
reg [10:0] m37_22;
reg [10:0] m37_23;
reg [10:0] m37_24;
reg [10:0] m38_0;
reg [10:0] m38_1;
reg [10:0] m38_2;
reg [10:0] m38_3;
reg [10:0] m38_4;
reg [10:0] m38_5;
reg [10:0] m38_6;
reg [10:0] m38_7;
reg [10:0] m38_8;
reg [10:0] m38_9;
reg [10:0] m38_10;
reg [10:0] m38_11;
reg [10:0] m38_12;
reg [10:0] m38_13;
reg [10:0] m38_14;
reg [10:0] m38_15;
reg [10:0] m38_16;
reg [10:0] m38_17;
reg [10:0] m38_18;
reg [10:0] m38_19;
reg [10:0] m38_20;
reg [10:0] m38_21;
reg [10:0] m38_22;
reg [10:0] m38_23;
reg [10:0] m38_24;
reg [10:0] m39_0;
reg [10:0] m39_1;
reg [10:0] m39_2;
reg [10:0] m39_3;
reg [10:0] m39_4;
reg [10:0] m39_5;
reg [10:0] m39_6;
reg [10:0] m39_7;
reg [10:0] m39_8;
reg [10:0] m39_9;
reg [10:0] m39_10;
reg [10:0] m39_11;
reg [10:0] m39_12;
reg [10:0] m39_13;
reg [10:0] m39_14;
reg [10:0] m39_15;
reg [10:0] m39_16;
reg [10:0] m39_17;
reg [10:0] m39_18;
reg [10:0] m39_19;
reg [10:0] m39_20;
reg [10:0] m39_21;
reg [10:0] m39_22;
reg [10:0] m39_23;
reg [10:0] m39_24;


 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_0<=891;io0[0:0]<=1;end
else if(m0_0<1250)begin m0_0<=m0_0+1;end
else if(m0_0==1250)begin m0_0<=0;io0[0:0]<=~io0[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_1<=1020;io0[1:1]<=0;end
else if(m0_1<1250)begin m0_1<=m0_1+1;end
else if(m0_1==1250)begin m0_1<=0;io0[1:1]<=~io0[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_2<=927;io0[2:2]<=1;end
else if(m0_2<1250)begin m0_2<=m0_2+1;end
else if(m0_2==1250)begin m0_2<=0;io0[2:2]<=~io0[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_3<=1225;io0[3:3]<=1;end
else if(m0_3<1250)begin m0_3<=m0_3+1;end
else if(m0_3==1250)begin m0_3<=0;io0[3:3]<=~io0[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_4<=1010;io0[4:4]<=1;end
else if(m0_4<1250)begin m0_4<=m0_4+1;end
else if(m0_4==1250)begin m0_4<=0;io0[4:4]<=~io0[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_5<=1138;io0[5:5]<=0;end
else if(m0_5<1250)begin m0_5<=m0_5+1;end
else if(m0_5==1250)begin m0_5<=0;io0[5:5]<=~io0[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_6<=12;io0[6:6]<=1;end
else if(m0_6<1250)begin m0_6<=m0_6+1;end
else if(m0_6==1250)begin m0_6<=0;io0[6:6]<=~io0[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_7<=624;io0[7:7]<=0;end
else if(m0_7<1250)begin m0_7<=m0_7+1;end
else if(m0_7==1250)begin m0_7<=0;io0[7:7]<=~io0[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_8<=992;io0[8:8]<=1;end
else if(m0_8<1250)begin m0_8<=m0_8+1;end
else if(m0_8==1250)begin m0_8<=0;io0[8:8]<=~io0[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_9<=959;io0[9:9]<=0;end
else if(m0_9<1250)begin m0_9<=m0_9+1;end
else if(m0_9==1250)begin m0_9<=0;io0[9:9]<=~io0[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_10<=246;io0[10:10]<=0;end
else if(m0_10<1250)begin m0_10<=m0_10+1;end
else if(m0_10==1250)begin m0_10<=0;io0[10:10]<=~io0[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_11<=322;io0[11:11]<=1;end
else if(m0_11<1250)begin m0_11<=m0_11+1;end
else if(m0_11==1250)begin m0_11<=0;io0[11:11]<=~io0[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_12<=103;io0[12:12]<=0;end
else if(m0_12<1250)begin m0_12<=m0_12+1;end
else if(m0_12==1250)begin m0_12<=0;io0[12:12]<=~io0[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_13<=260;io0[13:13]<=0;end
else if(m0_13<1250)begin m0_13<=m0_13+1;end
else if(m0_13==1250)begin m0_13<=0;io0[13:13]<=~io0[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_14<=215;io0[14:14]<=0;end
else if(m0_14<1250)begin m0_14<=m0_14+1;end
else if(m0_14==1250)begin m0_14<=0;io0[14:14]<=~io0[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_15<=419;io0[15:15]<=0;end
else if(m0_15<1250)begin m0_15<=m0_15+1;end
else if(m0_15==1250)begin m0_15<=0;io0[15:15]<=~io0[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_16<=762;io0[16:16]<=1;end
else if(m0_16<1250)begin m0_16<=m0_16+1;end
else if(m0_16==1250)begin m0_16<=0;io0[16:16]<=~io0[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_17<=90;io0[17:17]<=0;end
else if(m0_17<1250)begin m0_17<=m0_17+1;end
else if(m0_17==1250)begin m0_17<=0;io0[17:17]<=~io0[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_18<=442;io0[18:18]<=0;end
else if(m0_18<1250)begin m0_18<=m0_18+1;end
else if(m0_18==1250)begin m0_18<=0;io0[18:18]<=~io0[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_19<=297;io0[19:19]<=0;end
else if(m0_19<1250)begin m0_19<=m0_19+1;end
else if(m0_19==1250)begin m0_19<=0;io0[19:19]<=~io0[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_20<=377;io0[20:20]<=1;end
else if(m0_20<1250)begin m0_20<=m0_20+1;end
else if(m0_20==1250)begin m0_20<=0;io0[20:20]<=~io0[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_21<=420;io0[21:21]<=0;end
else if(m0_21<1250)begin m0_21<=m0_21+1;end
else if(m0_21==1250)begin m0_21<=0;io0[21:21]<=~io0[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_22<=1221;io0[22:22]<=0;end
else if(m0_22<1250)begin m0_22<=m0_22+1;end
else if(m0_22==1250)begin m0_22<=0;io0[22:22]<=~io0[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_23<=1238;io0[23:23]<=0;end
else if(m0_23<1250)begin m0_23<=m0_23+1;end
else if(m0_23==1250)begin m0_23<=0;io0[23:23]<=~io0[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m0_24<=99;io0[24:24]<=1;end
else if(m0_24<1250)begin m0_24<=m0_24+1;end
else if(m0_24==1250)begin m0_24<=0;io0[24:24]<=~io0[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_0<=984;io1[0:0]<=1;end
else if(m1_0<1250)begin m1_0<=m1_0+1;end
else if(m1_0==1250)begin m1_0<=0;io1[0:0]<=~io1[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_1<=1247;io1[1:1]<=0;end
else if(m1_1<1250)begin m1_1<=m1_1+1;end
else if(m1_1==1250)begin m1_1<=0;io1[1:1]<=~io1[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_2<=1171;io1[2:2]<=1;end
else if(m1_2<1250)begin m1_2<=m1_2+1;end
else if(m1_2==1250)begin m1_2<=0;io1[2:2]<=~io1[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_3<=308;io1[3:3]<=0;end
else if(m1_3<1250)begin m1_3<=m1_3+1;end
else if(m1_3==1250)begin m1_3<=0;io1[3:3]<=~io1[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_4<=142;io1[4:4]<=0;end
else if(m1_4<1250)begin m1_4<=m1_4+1;end
else if(m1_4==1250)begin m1_4<=0;io1[4:4]<=~io1[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_5<=300;io1[5:5]<=1;end
else if(m1_5<1250)begin m1_5<=m1_5+1;end
else if(m1_5==1250)begin m1_5<=0;io1[5:5]<=~io1[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_6<=346;io1[6:6]<=1;end
else if(m1_6<1250)begin m1_6<=m1_6+1;end
else if(m1_6==1250)begin m1_6<=0;io1[6:6]<=~io1[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_7<=895;io1[7:7]<=0;end
else if(m1_7<1250)begin m1_7<=m1_7+1;end
else if(m1_7==1250)begin m1_7<=0;io1[7:7]<=~io1[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_8<=1209;io1[8:8]<=1;end
else if(m1_8<1250)begin m1_8<=m1_8+1;end
else if(m1_8==1250)begin m1_8<=0;io1[8:8]<=~io1[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_9<=1143;io1[9:9]<=0;end
else if(m1_9<1250)begin m1_9<=m1_9+1;end
else if(m1_9==1250)begin m1_9<=0;io1[9:9]<=~io1[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_10<=641;io1[10:10]<=0;end
else if(m1_10<1250)begin m1_10<=m1_10+1;end
else if(m1_10==1250)begin m1_10<=0;io1[10:10]<=~io1[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_11<=679;io1[11:11]<=1;end
else if(m1_11<1250)begin m1_11<=m1_11+1;end
else if(m1_11==1250)begin m1_11<=0;io1[11:11]<=~io1[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_12<=383;io1[12:12]<=0;end
else if(m1_12<1250)begin m1_12<=m1_12+1;end
else if(m1_12==1250)begin m1_12<=0;io1[12:12]<=~io1[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_13<=452;io1[13:13]<=0;end
else if(m1_13<1250)begin m1_13<=m1_13+1;end
else if(m1_13==1250)begin m1_13<=0;io1[13:13]<=~io1[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_14<=382;io1[14:14]<=0;end
else if(m1_14<1250)begin m1_14<=m1_14+1;end
else if(m1_14==1250)begin m1_14<=0;io1[14:14]<=~io1[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_15<=816;io1[15:15]<=0;end
else if(m1_15<1250)begin m1_15<=m1_15+1;end
else if(m1_15==1250)begin m1_15<=0;io1[15:15]<=~io1[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_16<=1109;io1[16:16]<=1;end
else if(m1_16<1250)begin m1_16<=m1_16+1;end
else if(m1_16==1250)begin m1_16<=0;io1[16:16]<=~io1[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_17<=376;io1[17:17]<=0;end
else if(m1_17<1250)begin m1_17<=m1_17+1;end
else if(m1_17==1250)begin m1_17<=0;io1[17:17]<=~io1[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_18<=615;io1[18:18]<=0;end
else if(m1_18<1250)begin m1_18<=m1_18+1;end
else if(m1_18==1250)begin m1_18<=0;io1[18:18]<=~io1[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_19<=459;io1[19:19]<=0;end
else if(m1_19<1250)begin m1_19<=m1_19+1;end
else if(m1_19==1250)begin m1_19<=0;io1[19:19]<=~io1[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_20<=768;io1[20:20]<=1;end
else if(m1_20<1250)begin m1_20<=m1_20+1;end
else if(m1_20==1250)begin m1_20<=0;io1[20:20]<=~io1[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_21<=736;io1[21:21]<=0;end
else if(m1_21<1250)begin m1_21<=m1_21+1;end
else if(m1_21==1250)begin m1_21<=0;io1[21:21]<=~io1[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_22<=225;io1[22:22]<=1;end
else if(m1_22<1250)begin m1_22<=m1_22+1;end
else if(m1_22==1250)begin m1_22<=0;io1[22:22]<=~io1[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_23<=225;io1[23:23]<=1;end
else if(m1_23<1250)begin m1_23<=m1_23+1;end
else if(m1_23==1250)begin m1_23<=0;io1[23:23]<=~io1[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m1_24<=245;io1[24:24]<=1;end
else if(m1_24<1250)begin m1_24<=m1_24+1;end
else if(m1_24==1250)begin m1_24<=0;io1[24:24]<=~io1[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_0<=984;io2[0:0]<=1;end
else if(m2_0<1250)begin m2_0<=m2_0+1;end
else if(m2_0==1250)begin m2_0<=0;io2[0:0]<=~io2[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_1<=1247;io2[1:1]<=0;end
else if(m2_1<1250)begin m2_1<=m2_1+1;end
else if(m2_1==1250)begin m2_1<=0;io2[1:1]<=~io2[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_2<=1171;io2[2:2]<=1;end
else if(m2_2<1250)begin m2_2<=m2_2+1;end
else if(m2_2==1250)begin m2_2<=0;io2[2:2]<=~io2[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_3<=308;io2[3:3]<=0;end
else if(m2_3<1250)begin m2_3<=m2_3+1;end
else if(m2_3==1250)begin m2_3<=0;io2[3:3]<=~io2[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_4<=142;io2[4:4]<=0;end
else if(m2_4<1250)begin m2_4<=m2_4+1;end
else if(m2_4==1250)begin m2_4<=0;io2[4:4]<=~io2[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_5<=300;io2[5:5]<=1;end
else if(m2_5<1250)begin m2_5<=m2_5+1;end
else if(m2_5==1250)begin m2_5<=0;io2[5:5]<=~io2[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_6<=346;io2[6:6]<=1;end
else if(m2_6<1250)begin m2_6<=m2_6+1;end
else if(m2_6==1250)begin m2_6<=0;io2[6:6]<=~io2[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_7<=895;io2[7:7]<=0;end
else if(m2_7<1250)begin m2_7<=m2_7+1;end
else if(m2_7==1250)begin m2_7<=0;io2[7:7]<=~io2[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_8<=1209;io2[8:8]<=1;end
else if(m2_8<1250)begin m2_8<=m2_8+1;end
else if(m2_8==1250)begin m2_8<=0;io2[8:8]<=~io2[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_9<=1143;io2[9:9]<=0;end
else if(m2_9<1250)begin m2_9<=m2_9+1;end
else if(m2_9==1250)begin m2_9<=0;io2[9:9]<=~io2[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_10<=641;io2[10:10]<=0;end
else if(m2_10<1250)begin m2_10<=m2_10+1;end
else if(m2_10==1250)begin m2_10<=0;io2[10:10]<=~io2[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_11<=679;io2[11:11]<=1;end
else if(m2_11<1250)begin m2_11<=m2_11+1;end
else if(m2_11==1250)begin m2_11<=0;io2[11:11]<=~io2[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_12<=383;io2[12:12]<=0;end
else if(m2_12<1250)begin m2_12<=m2_12+1;end
else if(m2_12==1250)begin m2_12<=0;io2[12:12]<=~io2[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_13<=452;io2[13:13]<=0;end
else if(m2_13<1250)begin m2_13<=m2_13+1;end
else if(m2_13==1250)begin m2_13<=0;io2[13:13]<=~io2[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_14<=382;io2[14:14]<=0;end
else if(m2_14<1250)begin m2_14<=m2_14+1;end
else if(m2_14==1250)begin m2_14<=0;io2[14:14]<=~io2[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_15<=816;io2[15:15]<=0;end
else if(m2_15<1250)begin m2_15<=m2_15+1;end
else if(m2_15==1250)begin m2_15<=0;io2[15:15]<=~io2[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_16<=1109;io2[16:16]<=1;end
else if(m2_16<1250)begin m2_16<=m2_16+1;end
else if(m2_16==1250)begin m2_16<=0;io2[16:16]<=~io2[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_17<=376;io2[17:17]<=0;end
else if(m2_17<1250)begin m2_17<=m2_17+1;end
else if(m2_17==1250)begin m2_17<=0;io2[17:17]<=~io2[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_18<=615;io2[18:18]<=0;end
else if(m2_18<1250)begin m2_18<=m2_18+1;end
else if(m2_18==1250)begin m2_18<=0;io2[18:18]<=~io2[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_19<=459;io2[19:19]<=0;end
else if(m2_19<1250)begin m2_19<=m2_19+1;end
else if(m2_19==1250)begin m2_19<=0;io2[19:19]<=~io2[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_20<=768;io2[20:20]<=1;end
else if(m2_20<1250)begin m2_20<=m2_20+1;end
else if(m2_20==1250)begin m2_20<=0;io2[20:20]<=~io2[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_21<=736;io2[21:21]<=0;end
else if(m2_21<1250)begin m2_21<=m2_21+1;end
else if(m2_21==1250)begin m2_21<=0;io2[21:21]<=~io2[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_22<=225;io2[22:22]<=1;end
else if(m2_22<1250)begin m2_22<=m2_22+1;end
else if(m2_22==1250)begin m2_22<=0;io2[22:22]<=~io2[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_23<=225;io2[23:23]<=1;end
else if(m2_23<1250)begin m2_23<=m2_23+1;end
else if(m2_23==1250)begin m2_23<=0;io2[23:23]<=~io2[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m2_24<=245;io2[24:24]<=1;end
else if(m2_24<1250)begin m2_24<=m2_24+1;end
else if(m2_24==1250)begin m2_24<=0;io2[24:24]<=~io2[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_0<=893;io3[0:0]<=1;end
else if(m3_0<1250)begin m3_0<=m3_0+1;end
else if(m3_0==1250)begin m3_0<=0;io3[0:0]<=~io3[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_1<=1146;io3[1:1]<=0;end
else if(m3_1<1250)begin m3_1<=m3_1+1;end
else if(m3_1==1250)begin m3_1<=0;io3[1:1]<=~io3[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_2<=1073;io3[2:2]<=1;end
else if(m3_2<1250)begin m3_2<=m3_2+1;end
else if(m3_2==1250)begin m3_2<=0;io3[2:2]<=~io3[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_3<=388;io3[3:3]<=0;end
else if(m3_3<1250)begin m3_3<=m3_3+1;end
else if(m3_3==1250)begin m3_3<=0;io3[3:3]<=~io3[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_4<=177;io3[4:4]<=0;end
else if(m3_4<1250)begin m3_4<=m3_4+1;end
else if(m3_4==1250)begin m3_4<=0;io3[4:4]<=~io3[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_5<=445;io3[5:5]<=1;end
else if(m3_5<1250)begin m3_5<=m3_5+1;end
else if(m3_5==1250)begin m3_5<=0;io3[5:5]<=~io3[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_6<=391;io3[6:6]<=1;end
else if(m3_6<1250)begin m3_6<=m3_6+1;end
else if(m3_6==1250)begin m3_6<=0;io3[6:6]<=~io3[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_7<=910;io3[7:7]<=0;end
else if(m3_7<1250)begin m3_7<=m3_7+1;end
else if(m3_7==1250)begin m3_7<=0;io3[7:7]<=~io3[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_8<=1119;io3[8:8]<=1;end
else if(m3_8<1250)begin m3_8<=m3_8+1;end
else if(m3_8==1250)begin m3_8<=0;io3[8:8]<=~io3[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_9<=1099;io3[9:9]<=0;end
else if(m3_9<1250)begin m3_9<=m3_9+1;end
else if(m3_9==1250)begin m3_9<=0;io3[9:9]<=~io3[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_10<=844;io3[10:10]<=0;end
else if(m3_10<1250)begin m3_10<=m3_10+1;end
else if(m3_10==1250)begin m3_10<=0;io3[10:10]<=~io3[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_11<=812;io3[11:11]<=1;end
else if(m3_11<1250)begin m3_11<=m3_11+1;end
else if(m3_11==1250)begin m3_11<=0;io3[11:11]<=~io3[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_12<=428;io3[12:12]<=0;end
else if(m3_12<1250)begin m3_12<=m3_12+1;end
else if(m3_12==1250)begin m3_12<=0;io3[12:12]<=~io3[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_13<=420;io3[13:13]<=0;end
else if(m3_13<1250)begin m3_13<=m3_13+1;end
else if(m3_13==1250)begin m3_13<=0;io3[13:13]<=~io3[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_14<=251;io3[14:14]<=0;end
else if(m3_14<1250)begin m3_14<=m3_14+1;end
else if(m3_14==1250)begin m3_14<=0;io3[14:14]<=~io3[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_15<=1098;io3[15:15]<=0;end
else if(m3_15<1250)begin m3_15<=m3_15+1;end
else if(m3_15==1250)begin m3_15<=0;io3[15:15]<=~io3[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_16<=33;io3[16:16]<=0;end
else if(m3_16<1250)begin m3_16<=m3_16+1;end
else if(m3_16==1250)begin m3_16<=0;io3[16:16]<=~io3[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_17<=534;io3[17:17]<=0;end
else if(m3_17<1250)begin m3_17<=m3_17+1;end
else if(m3_17==1250)begin m3_17<=0;io3[17:17]<=~io3[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_18<=664;io3[18:18]<=0;end
else if(m3_18<1250)begin m3_18<=m3_18+1;end
else if(m3_18==1250)begin m3_18<=0;io3[18:18]<=~io3[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_19<=440;io3[19:19]<=0;end
else if(m3_19<1250)begin m3_19<=m3_19+1;end
else if(m3_19==1250)begin m3_19<=0;io3[19:19]<=~io3[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_20<=1035;io3[20:20]<=1;end
else if(m3_20<1250)begin m3_20<=m3_20+1;end
else if(m3_20==1250)begin m3_20<=0;io3[20:20]<=~io3[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_21<=966;io3[21:21]<=0;end
else if(m3_21<1250)begin m3_21<=m3_21+1;end
else if(m3_21==1250)begin m3_21<=0;io3[21:21]<=~io3[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_22<=379;io3[22:22]<=1;end
else if(m3_22<1250)begin m3_22<=m3_22+1;end
else if(m3_22==1250)begin m3_22<=0;io3[22:22]<=~io3[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_23<=368;io3[23:23]<=1;end
else if(m3_23<1250)begin m3_23<=m3_23+1;end
else if(m3_23==1250)begin m3_23<=0;io3[23:23]<=~io3[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m3_24<=296;io3[24:24]<=1;end
else if(m3_24<1250)begin m3_24<=m3_24+1;end
else if(m3_24==1250)begin m3_24<=0;io3[24:24]<=~io3[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_0<=597;io4[0:0]<=1;end
else if(m4_0<1250)begin m4_0<=m4_0+1;end
else if(m4_0==1250)begin m4_0<=0;io4[0:0]<=~io4[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_1<=833;io4[1:1]<=0;end
else if(m4_1<1250)begin m4_1<=m4_1+1;end
else if(m4_1==1250)begin m4_1<=0;io4[1:1]<=~io4[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_2<=788;io4[2:2]<=1;end
else if(m4_2<1250)begin m4_2<=m4_2+1;end
else if(m4_2==1250)begin m4_2<=0;io4[2:2]<=~io4[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_3<=252;io4[3:3]<=0;end
else if(m4_3<1250)begin m4_3<=m4_3+1;end
else if(m4_3==1250)begin m4_3<=0;io4[3:3]<=~io4[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_4<=12;io4[4:4]<=0;end
else if(m4_4<1250)begin m4_4<=m4_4+1;end
else if(m4_4==1250)begin m4_4<=0;io4[4:4]<=~io4[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_5<=294;io4[5:5]<=1;end
else if(m4_5<1250)begin m4_5<=m4_5+1;end
else if(m4_5==1250)begin m4_5<=0;io4[5:5]<=~io4[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_6<=158;io4[6:6]<=1;end
else if(m4_6<1250)begin m4_6<=m4_6+1;end
else if(m4_6==1250)begin m4_6<=0;io4[6:6]<=~io4[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_7<=658;io4[7:7]<=0;end
else if(m4_7<1250)begin m4_7<=m4_7+1;end
else if(m4_7==1250)begin m4_7<=0;io4[7:7]<=~io4[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_8<=793;io4[8:8]<=1;end
else if(m4_8<1250)begin m4_8<=m4_8+1;end
else if(m4_8==1250)begin m4_8<=0;io4[8:8]<=~io4[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_9<=724;io4[9:9]<=0;end
else if(m4_9<1250)begin m4_9<=m4_9+1;end
else if(m4_9==1250)begin m4_9<=0;io4[9:9]<=~io4[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_10<=719;io4[10:10]<=0;end
else if(m4_10<1250)begin m4_10<=m4_10+1;end
else if(m4_10==1250)begin m4_10<=0;io4[10:10]<=~io4[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_11<=622;io4[11:11]<=1;end
else if(m4_11<1250)begin m4_11<=m4_11+1;end
else if(m4_11==1250)begin m4_11<=0;io4[11:11]<=~io4[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_12<=184;io4[12:12]<=0;end
else if(m4_12<1250)begin m4_12<=m4_12+1;end
else if(m4_12==1250)begin m4_12<=0;io4[12:12]<=~io4[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_13<=101;io4[13:13]<=0;end
else if(m4_13<1250)begin m4_13<=m4_13+1;end
else if(m4_13==1250)begin m4_13<=0;io4[13:13]<=~io4[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_14<=1085;io4[14:14]<=1;end
else if(m4_14<1250)begin m4_14<=m4_14+1;end
else if(m4_14==1250)begin m4_14<=0;io4[14:14]<=~io4[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_15<=958;io4[15:15]<=0;end
else if(m4_15<1250)begin m4_15<=m4_15+1;end
else if(m4_15==1250)begin m4_15<=0;io4[15:15]<=~io4[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_16<=1076;io4[16:16]<=1;end
else if(m4_16<1250)begin m4_16<=m4_16+1;end
else if(m4_16==1250)begin m4_16<=0;io4[16:16]<=~io4[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_17<=301;io4[17:17]<=0;end
else if(m4_17<1250)begin m4_17<=m4_17+1;end
else if(m4_17==1250)begin m4_17<=0;io4[17:17]<=~io4[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_18<=341;io4[18:18]<=0;end
else if(m4_18<1250)begin m4_18<=m4_18+1;end
else if(m4_18==1250)begin m4_18<=0;io4[18:18]<=~io4[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_19<=24;io4[19:19]<=0;end
else if(m4_19<1250)begin m4_19<=m4_19+1;end
else if(m4_19==1250)begin m4_19<=0;io4[19:19]<=~io4[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_20<=857;io4[20:20]<=1;end
else if(m4_20<1250)begin m4_20<=m4_20+1;end
else if(m4_20==1250)begin m4_20<=0;io4[20:20]<=~io4[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_21<=748;io4[21:21]<=0;end
else if(m4_21<1250)begin m4_21<=m4_21+1;end
else if(m4_21==1250)begin m4_21<=0;io4[21:21]<=~io4[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_22<=107;io4[22:22]<=1;end
else if(m4_22<1250)begin m4_22<=m4_22+1;end
else if(m4_22==1250)begin m4_22<=0;io4[22:22]<=~io4[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_23<=48;io4[23:23]<=1;end
else if(m4_23<1250)begin m4_23<=m4_23+1;end
else if(m4_23==1250)begin m4_23<=0;io4[23:23]<=~io4[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m4_24<=1215;io4[24:24]<=0;end
else if(m4_24<1250)begin m4_24<=m4_24+1;end
else if(m4_24==1250)begin m4_24<=0;io4[24:24]<=~io4[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_0<=688;io5[0:0]<=1;end
else if(m5_0<1250)begin m5_0<=m5_0+1;end
else if(m5_0==1250)begin m5_0<=0;io5[0:0]<=~io5[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_1<=979;io5[1:1]<=0;end
else if(m5_1<1250)begin m5_1<=m5_1+1;end
else if(m5_1==1250)begin m5_1<=0;io5[1:1]<=~io5[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_2<=922;io5[2:2]<=1;end
else if(m5_2<1250)begin m5_2<=m5_2+1;end
else if(m5_2==1250)begin m5_2<=0;io5[2:2]<=~io5[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_3<=341;io5[3:3]<=0;end
else if(m5_3<1250)begin m5_3<=m5_3+1;end
else if(m5_3==1250)begin m5_3<=0;io5[3:3]<=~io5[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_4<=151;io5[4:4]<=0;end
else if(m5_4<1250)begin m5_4<=m5_4+1;end
else if(m5_4==1250)begin m5_4<=0;io5[4:4]<=~io5[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_5<=483;io5[5:5]<=1;end
else if(m5_5<1250)begin m5_5<=m5_5+1;end
else if(m5_5==1250)begin m5_5<=0;io5[5:5]<=~io5[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_6<=347;io5[6:6]<=1;end
else if(m5_6<1250)begin m5_6<=m5_6+1;end
else if(m5_6==1250)begin m5_6<=0;io5[6:6]<=~io5[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_7<=855;io5[7:7]<=0;end
else if(m5_7<1250)begin m5_7<=m5_7+1;end
else if(m5_7==1250)begin m5_7<=0;io5[7:7]<=~io5[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_8<=970;io5[8:8]<=1;end
else if(m5_8<1250)begin m5_8<=m5_8+1;end
else if(m5_8==1250)begin m5_8<=0;io5[8:8]<=~io5[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_9<=924;io5[9:9]<=0;end
else if(m5_9<1250)begin m5_9<=m5_9+1;end
else if(m5_9==1250)begin m5_9<=0;io5[9:9]<=~io5[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_10<=968;io5[10:10]<=0;end
else if(m5_10<1250)begin m5_10<=m5_10+1;end
else if(m5_10==1250)begin m5_10<=0;io5[10:10]<=~io5[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_11<=864;io5[11:11]<=1;end
else if(m5_11<1250)begin m5_11<=m5_11+1;end
else if(m5_11==1250)begin m5_11<=0;io5[11:11]<=~io5[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_12<=400;io5[12:12]<=0;end
else if(m5_12<1250)begin m5_12<=m5_12+1;end
else if(m5_12==1250)begin m5_12<=0;io5[12:12]<=~io5[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_13<=327;io5[13:13]<=0;end
else if(m5_13<1250)begin m5_13<=m5_13+1;end
else if(m5_13==1250)begin m5_13<=0;io5[13:13]<=~io5[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_14<=55;io5[14:14]<=0;end
else if(m5_14<1250)begin m5_14<=m5_14+1;end
else if(m5_14==1250)begin m5_14<=0;io5[14:14]<=~io5[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_15<=29;io5[15:15]<=1;end
else if(m5_15<1250)begin m5_15<=m5_15+1;end
else if(m5_15==1250)begin m5_15<=0;io5[15:15]<=~io5[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_16<=130;io5[16:16]<=0;end
else if(m5_16<1250)begin m5_16<=m5_16+1;end
else if(m5_16==1250)begin m5_16<=0;io5[16:16]<=~io5[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_17<=638;io5[17:17]<=0;end
else if(m5_17<1250)begin m5_17<=m5_17+1;end
else if(m5_17==1250)begin m5_17<=0;io5[17:17]<=~io5[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_18<=679;io5[18:18]<=0;end
else if(m5_18<1250)begin m5_18<=m5_18+1;end
else if(m5_18==1250)begin m5_18<=0;io5[18:18]<=~io5[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_19<=366;io5[19:19]<=0;end
else if(m5_19<1250)begin m5_19<=m5_19+1;end
else if(m5_19==1250)begin m5_19<=0;io5[19:19]<=~io5[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_20<=1223;io5[20:20]<=1;end
else if(m5_20<1250)begin m5_20<=m5_20+1;end
else if(m5_20==1250)begin m5_20<=0;io5[20:20]<=~io5[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_21<=1115;io5[21:21]<=0;end
else if(m5_21<1250)begin m5_21<=m5_21+1;end
else if(m5_21==1250)begin m5_21<=0;io5[21:21]<=~io5[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_22<=476;io5[22:22]<=1;end
else if(m5_22<1250)begin m5_22<=m5_22+1;end
else if(m5_22==1250)begin m5_22<=0;io5[22:22]<=~io5[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_23<=438;io5[23:23]<=1;end
else if(m5_23<1250)begin m5_23<=m5_23+1;end
else if(m5_23==1250)begin m5_23<=0;io5[23:23]<=~io5[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m5_24<=288;io5[24:24]<=1;end
else if(m5_24<1250)begin m5_24<=m5_24+1;end
else if(m5_24==1250)begin m5_24<=0;io5[24:24]<=~io5[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_0<=688;io6[0:0]<=1;end
else if(m6_0<1250)begin m6_0<=m6_0+1;end
else if(m6_0==1250)begin m6_0<=0;io6[0:0]<=~io6[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_1<=979;io6[1:1]<=0;end
else if(m6_1<1250)begin m6_1<=m6_1+1;end
else if(m6_1==1250)begin m6_1<=0;io6[1:1]<=~io6[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_2<=922;io6[2:2]<=1;end
else if(m6_2<1250)begin m6_2<=m6_2+1;end
else if(m6_2==1250)begin m6_2<=0;io6[2:2]<=~io6[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_3<=341;io6[3:3]<=0;end
else if(m6_3<1250)begin m6_3<=m6_3+1;end
else if(m6_3==1250)begin m6_3<=0;io6[3:3]<=~io6[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_4<=151;io6[4:4]<=0;end
else if(m6_4<1250)begin m6_4<=m6_4+1;end
else if(m6_4==1250)begin m6_4<=0;io6[4:4]<=~io6[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_5<=483;io6[5:5]<=1;end
else if(m6_5<1250)begin m6_5<=m6_5+1;end
else if(m6_5==1250)begin m6_5<=0;io6[5:5]<=~io6[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_6<=347;io6[6:6]<=1;end
else if(m6_6<1250)begin m6_6<=m6_6+1;end
else if(m6_6==1250)begin m6_6<=0;io6[6:6]<=~io6[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_7<=855;io6[7:7]<=0;end
else if(m6_7<1250)begin m6_7<=m6_7+1;end
else if(m6_7==1250)begin m6_7<=0;io6[7:7]<=~io6[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_8<=970;io6[8:8]<=1;end
else if(m6_8<1250)begin m6_8<=m6_8+1;end
else if(m6_8==1250)begin m6_8<=0;io6[8:8]<=~io6[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_9<=924;io6[9:9]<=0;end
else if(m6_9<1250)begin m6_9<=m6_9+1;end
else if(m6_9==1250)begin m6_9<=0;io6[9:9]<=~io6[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_10<=968;io6[10:10]<=0;end
else if(m6_10<1250)begin m6_10<=m6_10+1;end
else if(m6_10==1250)begin m6_10<=0;io6[10:10]<=~io6[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_11<=864;io6[11:11]<=1;end
else if(m6_11<1250)begin m6_11<=m6_11+1;end
else if(m6_11==1250)begin m6_11<=0;io6[11:11]<=~io6[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_12<=400;io6[12:12]<=0;end
else if(m6_12<1250)begin m6_12<=m6_12+1;end
else if(m6_12==1250)begin m6_12<=0;io6[12:12]<=~io6[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_13<=327;io6[13:13]<=0;end
else if(m6_13<1250)begin m6_13<=m6_13+1;end
else if(m6_13==1250)begin m6_13<=0;io6[13:13]<=~io6[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_14<=55;io6[14:14]<=0;end
else if(m6_14<1250)begin m6_14<=m6_14+1;end
else if(m6_14==1250)begin m6_14<=0;io6[14:14]<=~io6[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_15<=29;io6[15:15]<=1;end
else if(m6_15<1250)begin m6_15<=m6_15+1;end
else if(m6_15==1250)begin m6_15<=0;io6[15:15]<=~io6[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_16<=130;io6[16:16]<=0;end
else if(m6_16<1250)begin m6_16<=m6_16+1;end
else if(m6_16==1250)begin m6_16<=0;io6[16:16]<=~io6[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_17<=638;io6[17:17]<=0;end
else if(m6_17<1250)begin m6_17<=m6_17+1;end
else if(m6_17==1250)begin m6_17<=0;io6[17:17]<=~io6[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_18<=679;io6[18:18]<=0;end
else if(m6_18<1250)begin m6_18<=m6_18+1;end
else if(m6_18==1250)begin m6_18<=0;io6[18:18]<=~io6[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_19<=366;io6[19:19]<=0;end
else if(m6_19<1250)begin m6_19<=m6_19+1;end
else if(m6_19==1250)begin m6_19<=0;io6[19:19]<=~io6[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_20<=1223;io6[20:20]<=1;end
else if(m6_20<1250)begin m6_20<=m6_20+1;end
else if(m6_20==1250)begin m6_20<=0;io6[20:20]<=~io6[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_21<=1115;io6[21:21]<=0;end
else if(m6_21<1250)begin m6_21<=m6_21+1;end
else if(m6_21==1250)begin m6_21<=0;io6[21:21]<=~io6[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_22<=476;io6[22:22]<=1;end
else if(m6_22<1250)begin m6_22<=m6_22+1;end
else if(m6_22==1250)begin m6_22<=0;io6[22:22]<=~io6[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_23<=438;io6[23:23]<=1;end
else if(m6_23<1250)begin m6_23<=m6_23+1;end
else if(m6_23==1250)begin m6_23<=0;io6[23:23]<=~io6[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m6_24<=288;io6[24:24]<=1;end
else if(m6_24<1250)begin m6_24<=m6_24+1;end
else if(m6_24==1250)begin m6_24<=0;io6[24:24]<=~io6[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_0<=37;io7[0:0]<=1;end
else if(m7_0<1250)begin m7_0<=m7_0+1;end
else if(m7_0==1250)begin m7_0<=0;io7[0:0]<=~io7[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_1<=421;io7[1:1]<=0;end
else if(m7_1<1250)begin m7_1<=m7_1+1;end
else if(m7_1==1250)begin m7_1<=0;io7[1:1]<=~io7[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_2<=429;io7[2:2]<=1;end
else if(m7_2<1250)begin m7_2<=m7_2+1;end
else if(m7_2==1250)begin m7_2<=0;io7[2:2]<=~io7[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_3<=1109;io7[3:3]<=1;end
else if(m7_3<1250)begin m7_3<=m7_3+1;end
else if(m7_3==1250)begin m7_3<=0;io7[3:3]<=~io7[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_4<=1042;io7[4:4]<=1;end
else if(m7_4<1250)begin m7_4<=m7_4+1;end
else if(m7_4==1250)begin m7_4<=0;io7[4:4]<=~io7[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_5<=134;io7[5:5]<=1;end
else if(m7_5<1250)begin m7_5<=m7_5+1;end
else if(m7_5==1250)begin m7_5<=0;io7[5:5]<=~io7[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_6<=1197;io7[6:6]<=0;end
else if(m7_6<1250)begin m7_6<=m7_6+1;end
else if(m7_6==1250)begin m7_6<=0;io7[6:6]<=~io7[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_7<=430;io7[7:7]<=0;end
else if(m7_7<1250)begin m7_7<=m7_7+1;end
else if(m7_7==1250)begin m7_7<=0;io7[7:7]<=~io7[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_8<=492;io7[8:8]<=1;end
else if(m7_8<1250)begin m7_8<=m7_8+1;end
else if(m7_8==1250)begin m7_8<=0;io7[8:8]<=~io7[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_9<=286;io7[9:9]<=0;end
else if(m7_9<1250)begin m7_9<=m7_9+1;end
else if(m7_9==1250)begin m7_9<=0;io7[9:9]<=~io7[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_10<=703;io7[10:10]<=0;end
else if(m7_10<1250)begin m7_10<=m7_10+1;end
else if(m7_10==1250)begin m7_10<=0;io7[10:10]<=~io7[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_11<=562;io7[11:11]<=1;end
else if(m7_11<1250)begin m7_11<=m7_11+1;end
else if(m7_11==1250)begin m7_11<=0;io7[11:11]<=~io7[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_12<=24;io7[12:12]<=0;end
else if(m7_12<1250)begin m7_12<=m7_12+1;end
else if(m7_12==1250)begin m7_12<=0;io7[12:12]<=~io7[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_13<=1148;io7[13:13]<=1;end
else if(m7_13<1250)begin m7_13<=m7_13+1;end
else if(m7_13==1250)begin m7_13<=0;io7[13:13]<=~io7[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_14<=787;io7[14:14]<=1;end
else if(m7_14<1250)begin m7_14<=m7_14+1;end
else if(m7_14==1250)begin m7_14<=0;io7[14:14]<=~io7[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_15<=1054;io7[15:15]<=0;end
else if(m7_15<1250)begin m7_15<=m7_15+1;end
else if(m7_15==1250)begin m7_15<=0;io7[15:15]<=~io7[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_16<=1143;io7[16:16]<=1;end
else if(m7_16<1250)begin m7_16<=m7_16+1;end
else if(m7_16==1250)begin m7_16<=0;io7[16:16]<=~io7[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_17<=361;io7[17:17]<=0;end
else if(m7_17<1250)begin m7_17<=m7_17+1;end
else if(m7_17==1250)begin m7_17<=0;io7[17:17]<=~io7[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_18<=358;io7[18:18]<=0;end
else if(m7_18<1250)begin m7_18<=m7_18+1;end
else if(m7_18==1250)begin m7_18<=0;io7[18:18]<=~io7[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_19<=1200;io7[19:19]<=1;end
else if(m7_19<1250)begin m7_19<=m7_19+1;end
else if(m7_19==1250)begin m7_19<=0;io7[19:19]<=~io7[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_20<=1101;io7[20:20]<=1;end
else if(m7_20<1250)begin m7_20<=m7_20+1;end
else if(m7_20==1250)begin m7_20<=0;io7[20:20]<=~io7[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_21<=919;io7[21:21]<=0;end
else if(m7_21<1250)begin m7_21<=m7_21+1;end
else if(m7_21==1250)begin m7_21<=0;io7[21:21]<=~io7[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_22<=254;io7[22:22]<=1;end
else if(m7_22<1250)begin m7_22<=m7_22+1;end
else if(m7_22==1250)begin m7_22<=0;io7[22:22]<=~io7[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_23<=139;io7[23:23]<=1;end
else if(m7_23<1250)begin m7_23<=m7_23+1;end
else if(m7_23==1250)begin m7_23<=0;io7[23:23]<=~io7[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m7_24<=1196;io7[24:24]<=0;end
else if(m7_24<1250)begin m7_24<=m7_24+1;end
else if(m7_24==1250)begin m7_24<=0;io7[24:24]<=~io7[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_0<=37;io8[0:0]<=1;end
else if(m8_0<1250)begin m8_0<=m8_0+1;end
else if(m8_0==1250)begin m8_0<=0;io8[0:0]<=~io8[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_1<=421;io8[1:1]<=0;end
else if(m8_1<1250)begin m8_1<=m8_1+1;end
else if(m8_1==1250)begin m8_1<=0;io8[1:1]<=~io8[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_2<=429;io8[2:2]<=1;end
else if(m8_2<1250)begin m8_2<=m8_2+1;end
else if(m8_2==1250)begin m8_2<=0;io8[2:2]<=~io8[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_3<=1109;io8[3:3]<=1;end
else if(m8_3<1250)begin m8_3<=m8_3+1;end
else if(m8_3==1250)begin m8_3<=0;io8[3:3]<=~io8[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_4<=1042;io8[4:4]<=1;end
else if(m8_4<1250)begin m8_4<=m8_4+1;end
else if(m8_4==1250)begin m8_4<=0;io8[4:4]<=~io8[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_5<=134;io8[5:5]<=1;end
else if(m8_5<1250)begin m8_5<=m8_5+1;end
else if(m8_5==1250)begin m8_5<=0;io8[5:5]<=~io8[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_6<=1197;io8[6:6]<=0;end
else if(m8_6<1250)begin m8_6<=m8_6+1;end
else if(m8_6==1250)begin m8_6<=0;io8[6:6]<=~io8[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_7<=430;io8[7:7]<=0;end
else if(m8_7<1250)begin m8_7<=m8_7+1;end
else if(m8_7==1250)begin m8_7<=0;io8[7:7]<=~io8[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_8<=492;io8[8:8]<=1;end
else if(m8_8<1250)begin m8_8<=m8_8+1;end
else if(m8_8==1250)begin m8_8<=0;io8[8:8]<=~io8[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_9<=286;io8[9:9]<=0;end
else if(m8_9<1250)begin m8_9<=m8_9+1;end
else if(m8_9==1250)begin m8_9<=0;io8[9:9]<=~io8[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_10<=703;io8[10:10]<=0;end
else if(m8_10<1250)begin m8_10<=m8_10+1;end
else if(m8_10==1250)begin m8_10<=0;io8[10:10]<=~io8[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_11<=562;io8[11:11]<=1;end
else if(m8_11<1250)begin m8_11<=m8_11+1;end
else if(m8_11==1250)begin m8_11<=0;io8[11:11]<=~io8[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_12<=24;io8[12:12]<=0;end
else if(m8_12<1250)begin m8_12<=m8_12+1;end
else if(m8_12==1250)begin m8_12<=0;io8[12:12]<=~io8[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_13<=1148;io8[13:13]<=1;end
else if(m8_13<1250)begin m8_13<=m8_13+1;end
else if(m8_13==1250)begin m8_13<=0;io8[13:13]<=~io8[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_14<=787;io8[14:14]<=1;end
else if(m8_14<1250)begin m8_14<=m8_14+1;end
else if(m8_14==1250)begin m8_14<=0;io8[14:14]<=~io8[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_15<=1054;io8[15:15]<=0;end
else if(m8_15<1250)begin m8_15<=m8_15+1;end
else if(m8_15==1250)begin m8_15<=0;io8[15:15]<=~io8[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_16<=1143;io8[16:16]<=1;end
else if(m8_16<1250)begin m8_16<=m8_16+1;end
else if(m8_16==1250)begin m8_16<=0;io8[16:16]<=~io8[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_17<=361;io8[17:17]<=0;end
else if(m8_17<1250)begin m8_17<=m8_17+1;end
else if(m8_17==1250)begin m8_17<=0;io8[17:17]<=~io8[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_18<=358;io8[18:18]<=0;end
else if(m8_18<1250)begin m8_18<=m8_18+1;end
else if(m8_18==1250)begin m8_18<=0;io8[18:18]<=~io8[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_19<=1200;io8[19:19]<=1;end
else if(m8_19<1250)begin m8_19<=m8_19+1;end
else if(m8_19==1250)begin m8_19<=0;io8[19:19]<=~io8[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_20<=1101;io8[20:20]<=1;end
else if(m8_20<1250)begin m8_20<=m8_20+1;end
else if(m8_20==1250)begin m8_20<=0;io8[20:20]<=~io8[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_21<=919;io8[21:21]<=0;end
else if(m8_21<1250)begin m8_21<=m8_21+1;end
else if(m8_21==1250)begin m8_21<=0;io8[21:21]<=~io8[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_22<=254;io8[22:22]<=1;end
else if(m8_22<1250)begin m8_22<=m8_22+1;end
else if(m8_22==1250)begin m8_22<=0;io8[22:22]<=~io8[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_23<=139;io8[23:23]<=1;end
else if(m8_23<1250)begin m8_23<=m8_23+1;end
else if(m8_23==1250)begin m8_23<=0;io8[23:23]<=~io8[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m8_24<=1196;io8[24:24]<=0;end
else if(m8_24<1250)begin m8_24<=m8_24+1;end
else if(m8_24==1250)begin m8_24<=0;io8[24:24]<=~io8[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_0<=1106;io9[0:0]<=0;end
else if(m9_0<1250)begin m9_0<=m9_0+1;end
else if(m9_0==1250)begin m9_0<=0;io9[0:0]<=~io9[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_1<=277;io9[1:1]<=0;end
else if(m9_1<1250)begin m9_1<=m9_1+1;end
else if(m9_1==1250)begin m9_1<=0;io9[1:1]<=~io9[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_2<=282;io9[2:2]<=1;end
else if(m9_2<1250)begin m9_2<=m9_2+1;end
else if(m9_2==1250)begin m9_2<=0;io9[2:2]<=~io9[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_3<=940;io9[3:3]<=1;end
else if(m9_3<1250)begin m9_3<=m9_3+1;end
else if(m9_3==1250)begin m9_3<=0;io9[3:3]<=~io9[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_4<=920;io9[4:4]<=1;end
else if(m9_4<1250)begin m9_4<=m9_4+1;end
else if(m9_4==1250)begin m9_4<=0;io9[4:4]<=~io9[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_5<=75;io9[5:5]<=1;end
else if(m9_5<1250)begin m9_5<=m9_5+1;end
else if(m9_5==1250)begin m9_5<=0;io9[5:5]<=~io9[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_6<=1102;io9[6:6]<=0;end
else if(m9_6<1250)begin m9_6<=m9_6+1;end
else if(m9_6==1250)begin m9_6<=0;io9[6:6]<=~io9[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_7<=361;io9[7:7]<=0;end
else if(m9_7<1250)begin m9_7<=m9_7+1;end
else if(m9_7==1250)begin m9_7<=0;io9[7:7]<=~io9[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_8<=420;io9[8:8]<=1;end
else if(m9_8<1250)begin m9_8<=m9_8+1;end
else if(m9_8==1250)begin m9_8<=0;io9[8:8]<=~io9[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_9<=158;io9[9:9]<=0;end
else if(m9_9<1250)begin m9_9<=m9_9+1;end
else if(m9_9==1250)begin m9_9<=0;io9[9:9]<=~io9[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_10<=703;io9[10:10]<=0;end
else if(m9_10<1250)begin m9_10<=m9_10+1;end
else if(m9_10==1250)begin m9_10<=0;io9[10:10]<=~io9[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_11<=562;io9[11:11]<=1;end
else if(m9_11<1250)begin m9_11<=m9_11+1;end
else if(m9_11==1250)begin m9_11<=0;io9[11:11]<=~io9[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_12<=24;io9[12:12]<=0;end
else if(m9_12<1250)begin m9_12<=m9_12+1;end
else if(m9_12==1250)begin m9_12<=0;io9[12:12]<=~io9[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_13<=1148;io9[13:13]<=1;end
else if(m9_13<1250)begin m9_13<=m9_13+1;end
else if(m9_13==1250)begin m9_13<=0;io9[13:13]<=~io9[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_14<=787;io9[14:14]<=1;end
else if(m9_14<1250)begin m9_14<=m9_14+1;end
else if(m9_14==1250)begin m9_14<=0;io9[14:14]<=~io9[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_15<=1113;io9[15:15]<=0;end
else if(m9_15<1250)begin m9_15<=m9_15+1;end
else if(m9_15==1250)begin m9_15<=0;io9[15:15]<=~io9[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_16<=1238;io9[16:16]<=1;end
else if(m9_16<1250)begin m9_16<=m9_16+1;end
else if(m9_16==1250)begin m9_16<=0;io9[16:16]<=~io9[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_17<=430;io9[17:17]<=0;end
else if(m9_17<1250)begin m9_17<=m9_17+1;end
else if(m9_17==1250)begin m9_17<=0;io9[17:17]<=~io9[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_18<=430;io9[18:18]<=0;end
else if(m9_18<1250)begin m9_18<=m9_18+1;end
else if(m9_18==1250)begin m9_18<=0;io9[18:18]<=~io9[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_19<=77;io9[19:19]<=0;end
else if(m9_19<1250)begin m9_19<=m9_19+1;end
else if(m9_19==1250)begin m9_19<=0;io9[19:19]<=~io9[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_20<=1222;io9[20:20]<=1;end
else if(m9_20<1250)begin m9_20<=m9_20+1;end
else if(m9_20==1250)begin m9_20<=0;io9[20:20]<=~io9[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_21<=1088;io9[21:21]<=0;end
else if(m9_21<1250)begin m9_21<=m9_21+1;end
else if(m9_21==1250)begin m9_21<=0;io9[21:21]<=~io9[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_22<=401;io9[22:22]<=1;end
else if(m9_22<1250)begin m9_22<=m9_22+1;end
else if(m9_22==1250)begin m9_22<=0;io9[22:22]<=~io9[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_23<=282;io9[23:23]<=1;end
else if(m9_23<1250)begin m9_23<=m9_23+1;end
else if(m9_23==1250)begin m9_23<=0;io9[23:23]<=~io9[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m9_24<=127;io9[24:24]<=1;end
else if(m9_24<1250)begin m9_24<=m9_24+1;end
else if(m9_24==1250)begin m9_24<=0;io9[24:24]<=~io9[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_0<=888;io10[0:0]<=0;end
else if(m10_0<1250)begin m10_0<=m10_0+1;end
else if(m10_0==1250)begin m10_0<=0;io10[0:0]<=~io10[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_1<=14;io10[1:1]<=0;end
else if(m10_1<1250)begin m10_1<=m10_1+1;end
else if(m10_1==1250)begin m10_1<=0;io10[1:1]<=~io10[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_2<=28;io10[2:2]<=1;end
else if(m10_2<1250)begin m10_2<=m10_2+1;end
else if(m10_2==1250)begin m10_2<=0;io10[2:2]<=~io10[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_3<=712;io10[3:3]<=1;end
else if(m10_3<1250)begin m10_3<=m10_3+1;end
else if(m10_3==1250)begin m10_3<=0;io10[3:3]<=~io10[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_4<=677;io10[4:4]<=1;end
else if(m10_4<1250)begin m10_4<=m10_4+1;end
else if(m10_4==1250)begin m10_4<=0;io10[4:4]<=~io10[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_5<=1155;io10[5:5]<=0;end
else if(m10_5<1250)begin m10_5<=m10_5+1;end
else if(m10_5==1250)begin m10_5<=0;io10[5:5]<=~io10[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_6<=911;io10[6:6]<=0;end
else if(m10_6<1250)begin m10_6<=m10_6+1;end
else if(m10_6==1250)begin m10_6<=0;io10[6:6]<=~io10[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_7<=168;io10[7:7]<=0;end
else if(m10_7<1250)begin m10_7<=m10_7+1;end
else if(m10_7==1250)begin m10_7<=0;io10[7:7]<=~io10[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_8<=227;io10[8:8]<=1;end
else if(m10_8<1250)begin m10_8<=m10_8+1;end
else if(m10_8==1250)begin m10_8<=0;io10[8:8]<=~io10[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_9<=1185;io10[9:9]<=1;end
else if(m10_9<1250)begin m10_9<=m10_9+1;end
else if(m10_9==1250)begin m10_9<=0;io10[9:9]<=~io10[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_10<=597;io10[10:10]<=0;end
else if(m10_10<1250)begin m10_10<=m10_10+1;end
else if(m10_10==1250)begin m10_10<=0;io10[10:10]<=~io10[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_11<=453;io10[11:11]<=1;end
else if(m10_11<1250)begin m10_11<=m10_11+1;end
else if(m10_11==1250)begin m10_11<=0;io10[11:11]<=~io10[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_12<=1183;io10[12:12]<=1;end
else if(m10_12<1250)begin m10_12<=m10_12+1;end
else if(m10_12==1250)begin m10_12<=0;io10[12:12]<=~io10[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_13<=1054;io10[13:13]<=1;end
else if(m10_13<1250)begin m10_13<=m10_13+1;end
else if(m10_13==1250)begin m10_13<=0;io10[13:13]<=~io10[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_14<=682;io10[14:14]<=1;end
else if(m10_14<1250)begin m10_14<=m10_14+1;end
else if(m10_14==1250)begin m10_14<=0;io10[14:14]<=~io10[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_15<=1066;io10[15:15]<=0;end
else if(m10_15<1250)begin m10_15<=m10_15+1;end
else if(m10_15==1250)begin m10_15<=0;io10[15:15]<=~io10[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_16<=1212;io10[16:16]<=1;end
else if(m10_16<1250)begin m10_16<=m10_16+1;end
else if(m10_16==1250)begin m10_16<=0;io10[16:16]<=~io10[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_17<=377;io10[17:17]<=0;end
else if(m10_17<1250)begin m10_17<=m10_17+1;end
else if(m10_17==1250)begin m10_17<=0;io10[17:17]<=~io10[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_18<=383;io10[18:18]<=0;end
else if(m10_18<1250)begin m10_18<=m10_18+1;end
else if(m10_18==1250)begin m10_18<=0;io10[18:18]<=~io10[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_19<=67;io10[19:19]<=0;end
else if(m10_19<1250)begin m10_19<=m10_19+1;end
else if(m10_19==1250)begin m10_19<=0;io10[19:19]<=~io10[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_20<=1220;io10[20:20]<=1;end
else if(m10_20<1250)begin m10_20<=m10_20+1;end
else if(m10_20==1250)begin m10_20<=0;io10[20:20]<=~io10[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_21<=1204;io10[21:21]<=0;end
else if(m10_21<1250)begin m10_21<=m10_21+1;end
else if(m10_21==1250)begin m10_21<=0;io10[21:21]<=~io10[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_22<=419;io10[22:22]<=1;end
else if(m10_22<1250)begin m10_22<=m10_22+1;end
else if(m10_22==1250)begin m10_22<=0;io10[22:22]<=~io10[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_23<=290;io10[23:23]<=1;end
else if(m10_23<1250)begin m10_23<=m10_23+1;end
else if(m10_23==1250)begin m10_23<=0;io10[23:23]<=~io10[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m10_24<=254;io10[24:24]<=1;end
else if(m10_24<1250)begin m10_24<=m10_24+1;end
else if(m10_24==1250)begin m10_24<=0;io10[24:24]<=~io10[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_0<=888;io11[0:0]<=0;end
else if(m11_0<1250)begin m11_0<=m11_0+1;end
else if(m11_0==1250)begin m11_0<=0;io11[0:0]<=~io11[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_1<=14;io11[1:1]<=0;end
else if(m11_1<1250)begin m11_1<=m11_1+1;end
else if(m11_1==1250)begin m11_1<=0;io11[1:1]<=~io11[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_2<=28;io11[2:2]<=1;end
else if(m11_2<1250)begin m11_2<=m11_2+1;end
else if(m11_2==1250)begin m11_2<=0;io11[2:2]<=~io11[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_3<=712;io11[3:3]<=1;end
else if(m11_3<1250)begin m11_3<=m11_3+1;end
else if(m11_3==1250)begin m11_3<=0;io11[3:3]<=~io11[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_4<=677;io11[4:4]<=1;end
else if(m11_4<1250)begin m11_4<=m11_4+1;end
else if(m11_4==1250)begin m11_4<=0;io11[4:4]<=~io11[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_5<=1155;io11[5:5]<=0;end
else if(m11_5<1250)begin m11_5<=m11_5+1;end
else if(m11_5==1250)begin m11_5<=0;io11[5:5]<=~io11[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_6<=911;io11[6:6]<=0;end
else if(m11_6<1250)begin m11_6<=m11_6+1;end
else if(m11_6==1250)begin m11_6<=0;io11[6:6]<=~io11[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_7<=168;io11[7:7]<=0;end
else if(m11_7<1250)begin m11_7<=m11_7+1;end
else if(m11_7==1250)begin m11_7<=0;io11[7:7]<=~io11[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_8<=227;io11[8:8]<=1;end
else if(m11_8<1250)begin m11_8<=m11_8+1;end
else if(m11_8==1250)begin m11_8<=0;io11[8:8]<=~io11[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_9<=1185;io11[9:9]<=1;end
else if(m11_9<1250)begin m11_9<=m11_9+1;end
else if(m11_9==1250)begin m11_9<=0;io11[9:9]<=~io11[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_10<=597;io11[10:10]<=0;end
else if(m11_10<1250)begin m11_10<=m11_10+1;end
else if(m11_10==1250)begin m11_10<=0;io11[10:10]<=~io11[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_11<=453;io11[11:11]<=1;end
else if(m11_11<1250)begin m11_11<=m11_11+1;end
else if(m11_11==1250)begin m11_11<=0;io11[11:11]<=~io11[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_12<=1183;io11[12:12]<=1;end
else if(m11_12<1250)begin m11_12<=m11_12+1;end
else if(m11_12==1250)begin m11_12<=0;io11[12:12]<=~io11[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_13<=1054;io11[13:13]<=1;end
else if(m11_13<1250)begin m11_13<=m11_13+1;end
else if(m11_13==1250)begin m11_13<=0;io11[13:13]<=~io11[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_14<=682;io11[14:14]<=1;end
else if(m11_14<1250)begin m11_14<=m11_14+1;end
else if(m11_14==1250)begin m11_14<=0;io11[14:14]<=~io11[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_15<=1066;io11[15:15]<=0;end
else if(m11_15<1250)begin m11_15<=m11_15+1;end
else if(m11_15==1250)begin m11_15<=0;io11[15:15]<=~io11[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_16<=1212;io11[16:16]<=1;end
else if(m11_16<1250)begin m11_16<=m11_16+1;end
else if(m11_16==1250)begin m11_16<=0;io11[16:16]<=~io11[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_17<=377;io11[17:17]<=0;end
else if(m11_17<1250)begin m11_17<=m11_17+1;end
else if(m11_17==1250)begin m11_17<=0;io11[17:17]<=~io11[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_18<=383;io11[18:18]<=0;end
else if(m11_18<1250)begin m11_18<=m11_18+1;end
else if(m11_18==1250)begin m11_18<=0;io11[18:18]<=~io11[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_19<=67;io11[19:19]<=0;end
else if(m11_19<1250)begin m11_19<=m11_19+1;end
else if(m11_19==1250)begin m11_19<=0;io11[19:19]<=~io11[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_20<=1220;io11[20:20]<=1;end
else if(m11_20<1250)begin m11_20<=m11_20+1;end
else if(m11_20==1250)begin m11_20<=0;io11[20:20]<=~io11[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_21<=1204;io11[21:21]<=0;end
else if(m11_21<1250)begin m11_21<=m11_21+1;end
else if(m11_21==1250)begin m11_21<=0;io11[21:21]<=~io11[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_22<=419;io11[22:22]<=1;end
else if(m11_22<1250)begin m11_22<=m11_22+1;end
else if(m11_22==1250)begin m11_22<=0;io11[22:22]<=~io11[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_23<=290;io11[23:23]<=1;end
else if(m11_23<1250)begin m11_23<=m11_23+1;end
else if(m11_23==1250)begin m11_23<=0;io11[23:23]<=~io11[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m11_24<=254;io11[24:24]<=1;end
else if(m11_24<1250)begin m11_24<=m11_24+1;end
else if(m11_24==1250)begin m11_24<=0;io11[24:24]<=~io11[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_0<=1125;io12[0:0]<=0;end
else if(m12_0<1250)begin m12_0<=m12_0+1;end
else if(m12_0==1250)begin m12_0<=0;io12[0:0]<=~io12[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_1<=187;io12[1:1]<=0;end
else if(m12_1<1250)begin m12_1<=m12_1+1;end
else if(m12_1==1250)begin m12_1<=0;io12[1:1]<=~io12[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_2<=135;io12[2:2]<=1;end
else if(m12_2<1250)begin m12_2<=m12_2+1;end
else if(m12_2==1250)begin m12_2<=0;io12[2:2]<=~io12[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_3<=769;io12[3:3]<=1;end
else if(m12_3<1250)begin m12_3<=m12_3+1;end
else if(m12_3==1250)begin m12_3<=0;io12[3:3]<=~io12[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_4<=677;io12[4:4]<=1;end
else if(m12_4<1250)begin m12_4<=m12_4+1;end
else if(m12_4==1250)begin m12_4<=0;io12[4:4]<=~io12[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_5<=1229;io12[5:5]<=0;end
else if(m12_5<1250)begin m12_5<=m12_5+1;end
else if(m12_5==1250)begin m12_5<=0;io12[5:5]<=~io12[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_6<=1034;io12[6:6]<=0;end
else if(m12_6<1250)begin m12_6<=m12_6+1;end
else if(m12_6==1250)begin m12_6<=0;io12[6:6]<=~io12[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_7<=301;io12[7:7]<=0;end
else if(m12_7<1250)begin m12_7<=m12_7+1;end
else if(m12_7==1250)begin m12_7<=0;io12[7:7]<=~io12[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_8<=404;io12[8:8]<=1;end
else if(m12_8<1250)begin m12_8<=m12_8+1;end
else if(m12_8==1250)begin m12_8<=0;io12[8:8]<=~io12[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_9<=232;io12[9:9]<=0;end
else if(m12_9<1250)begin m12_9<=m12_9+1;end
else if(m12_9==1250)begin m12_9<=0;io12[9:9]<=~io12[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_10<=719;io12[10:10]<=0;end
else if(m12_10<1250)begin m12_10<=m12_10+1;end
else if(m12_10==1250)begin m12_10<=0;io12[10:10]<=~io12[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_11<=622;io12[11:11]<=1;end
else if(m12_11<1250)begin m12_11<=m12_11+1;end
else if(m12_11==1250)begin m12_11<=0;io12[11:11]<=~io12[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_12<=184;io12[12:12]<=0;end
else if(m12_12<1250)begin m12_12<=m12_12+1;end
else if(m12_12==1250)begin m12_12<=0;io12[12:12]<=~io12[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_13<=101;io12[13:13]<=0;end
else if(m12_13<1250)begin m12_13<=m12_13+1;end
else if(m12_13==1250)begin m12_13<=0;io12[13:13]<=~io12[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_14<=1085;io12[14:14]<=1;end
else if(m12_14<1250)begin m12_14<=m12_14+1;end
else if(m12_14==1250)begin m12_14<=0;io12[14:14]<=~io12[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_15<=23;io12[15:15]<=1;end
else if(m12_15<1250)begin m12_15<=m12_15+1;end
else if(m12_15==1250)begin m12_15<=0;io12[15:15]<=~io12[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_16<=200;io12[16:16]<=0;end
else if(m12_16<1250)begin m12_16<=m12_16+1;end
else if(m12_16==1250)begin m12_16<=0;io12[16:16]<=~io12[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_17<=658;io12[17:17]<=0;end
else if(m12_17<1250)begin m12_17<=m12_17+1;end
else if(m12_17==1250)begin m12_17<=0;io12[17:17]<=~io12[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_18<=731;io12[18:18]<=0;end
else if(m12_18<1250)begin m12_18<=m12_18+1;end
else if(m12_18==1250)begin m12_18<=0;io12[18:18]<=~io12[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_19<=516;io12[19:19]<=0;end
else if(m12_19<1250)begin m12_19<=m12_19+1;end
else if(m12_19==1250)begin m12_19<=0;io12[19:19]<=~io12[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_20<=192;io12[20:20]<=0;end
else if(m12_20<1250)begin m12_20<=m12_20+1;end
else if(m12_20==1250)begin m12_20<=0;io12[20:20]<=~io12[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_21<=231;io12[21:21]<=1;end
else if(m12_21<1250)begin m12_21<=m12_21+1;end
else if(m12_21==1250)begin m12_21<=0;io12[21:21]<=~io12[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_22<=760;io12[22:22]<=1;end
else if(m12_22<1250)begin m12_22<=m12_22+1;end
else if(m12_22==1250)begin m12_22<=0;io12[22:22]<=~io12[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_23<=695;io12[23:23]<=1;end
else if(m12_23<1250)begin m12_23<=m12_23+1;end
else if(m12_23==1250)begin m12_23<=0;io12[23:23]<=~io12[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m12_24<=687;io12[24:24]<=1;end
else if(m12_24<1250)begin m12_24<=m12_24+1;end
else if(m12_24==1250)begin m12_24<=0;io12[24:24]<=~io12[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_0<=1125;io13[0:0]<=0;end
else if(m13_0<1250)begin m13_0<=m13_0+1;end
else if(m13_0==1250)begin m13_0<=0;io13[0:0]<=~io13[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_1<=187;io13[1:1]<=0;end
else if(m13_1<1250)begin m13_1<=m13_1+1;end
else if(m13_1==1250)begin m13_1<=0;io13[1:1]<=~io13[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_2<=135;io13[2:2]<=1;end
else if(m13_2<1250)begin m13_2<=m13_2+1;end
else if(m13_2==1250)begin m13_2<=0;io13[2:2]<=~io13[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_3<=769;io13[3:3]<=1;end
else if(m13_3<1250)begin m13_3<=m13_3+1;end
else if(m13_3==1250)begin m13_3<=0;io13[3:3]<=~io13[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_4<=677;io13[4:4]<=1;end
else if(m13_4<1250)begin m13_4<=m13_4+1;end
else if(m13_4==1250)begin m13_4<=0;io13[4:4]<=~io13[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_5<=1229;io13[5:5]<=0;end
else if(m13_5<1250)begin m13_5<=m13_5+1;end
else if(m13_5==1250)begin m13_5<=0;io13[5:5]<=~io13[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_6<=1034;io13[6:6]<=0;end
else if(m13_6<1250)begin m13_6<=m13_6+1;end
else if(m13_6==1250)begin m13_6<=0;io13[6:6]<=~io13[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_7<=301;io13[7:7]<=0;end
else if(m13_7<1250)begin m13_7<=m13_7+1;end
else if(m13_7==1250)begin m13_7<=0;io13[7:7]<=~io13[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_8<=404;io13[8:8]<=1;end
else if(m13_8<1250)begin m13_8<=m13_8+1;end
else if(m13_8==1250)begin m13_8<=0;io13[8:8]<=~io13[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_9<=232;io13[9:9]<=0;end
else if(m13_9<1250)begin m13_9<=m13_9+1;end
else if(m13_9==1250)begin m13_9<=0;io13[9:9]<=~io13[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_10<=719;io13[10:10]<=0;end
else if(m13_10<1250)begin m13_10<=m13_10+1;end
else if(m13_10==1250)begin m13_10<=0;io13[10:10]<=~io13[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_11<=622;io13[11:11]<=1;end
else if(m13_11<1250)begin m13_11<=m13_11+1;end
else if(m13_11==1250)begin m13_11<=0;io13[11:11]<=~io13[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_12<=184;io13[12:12]<=0;end
else if(m13_12<1250)begin m13_12<=m13_12+1;end
else if(m13_12==1250)begin m13_12<=0;io13[12:12]<=~io13[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_13<=101;io13[13:13]<=0;end
else if(m13_13<1250)begin m13_13<=m13_13+1;end
else if(m13_13==1250)begin m13_13<=0;io13[13:13]<=~io13[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_14<=1085;io13[14:14]<=1;end
else if(m13_14<1250)begin m13_14<=m13_14+1;end
else if(m13_14==1250)begin m13_14<=0;io13[14:14]<=~io13[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_15<=23;io13[15:15]<=1;end
else if(m13_15<1250)begin m13_15<=m13_15+1;end
else if(m13_15==1250)begin m13_15<=0;io13[15:15]<=~io13[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_16<=200;io13[16:16]<=0;end
else if(m13_16<1250)begin m13_16<=m13_16+1;end
else if(m13_16==1250)begin m13_16<=0;io13[16:16]<=~io13[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_17<=658;io13[17:17]<=0;end
else if(m13_17<1250)begin m13_17<=m13_17+1;end
else if(m13_17==1250)begin m13_17<=0;io13[17:17]<=~io13[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_18<=731;io13[18:18]<=0;end
else if(m13_18<1250)begin m13_18<=m13_18+1;end
else if(m13_18==1250)begin m13_18<=0;io13[18:18]<=~io13[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_19<=516;io13[19:19]<=0;end
else if(m13_19<1250)begin m13_19<=m13_19+1;end
else if(m13_19==1250)begin m13_19<=0;io13[19:19]<=~io13[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_20<=192;io13[20:20]<=0;end
else if(m13_20<1250)begin m13_20<=m13_20+1;end
else if(m13_20==1250)begin m13_20<=0;io13[20:20]<=~io13[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_21<=231;io13[21:21]<=1;end
else if(m13_21<1250)begin m13_21<=m13_21+1;end
else if(m13_21==1250)begin m13_21<=0;io13[21:21]<=~io13[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_22<=760;io13[22:22]<=1;end
else if(m13_22<1250)begin m13_22<=m13_22+1;end
else if(m13_22==1250)begin m13_22<=0;io13[22:22]<=~io13[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_23<=695;io13[23:23]<=1;end
else if(m13_23<1250)begin m13_23<=m13_23+1;end
else if(m13_23==1250)begin m13_23<=0;io13[23:23]<=~io13[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m13_24<=687;io13[24:24]<=1;end
else if(m13_24<1250)begin m13_24<=m13_24+1;end
else if(m13_24==1250)begin m13_24<=0;io13[24:24]<=~io13[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_0<=1000;io14[0:0]<=0;end
else if(m14_0<1250)begin m14_0<=m14_0+1;end
else if(m14_0==1250)begin m14_0<=0;io14[0:0]<=~io14[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_1<=23;io14[1:1]<=0;end
else if(m14_1<1250)begin m14_1<=m14_1+1;end
else if(m14_1==1250)begin m14_1<=0;io14[1:1]<=~io14[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_2<=1231;io14[2:2]<=0;end
else if(m14_2<1250)begin m14_2<=m14_2+1;end
else if(m14_2==1250)begin m14_2<=0;io14[2:2]<=~io14[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_3<=576;io14[3:3]<=1;end
else if(m14_3<1250)begin m14_3<=m14_3+1;end
else if(m14_3==1250)begin m14_3<=0;io14[3:3]<=~io14[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_4<=520;io14[4:4]<=1;end
else if(m14_4<1250)begin m14_4<=m14_4+1;end
else if(m14_4==1250)begin m14_4<=0;io14[4:4]<=~io14[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_5<=1103;io14[5:5]<=0;end
else if(m14_5<1250)begin m14_5<=m14_5+1;end
else if(m14_5==1250)begin m14_5<=0;io14[5:5]<=~io14[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_6<=938;io14[6:6]<=0;end
else if(m14_6<1250)begin m14_6<=m14_6+1;end
else if(m14_6==1250)begin m14_6<=0;io14[6:6]<=~io14[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_7<=176;io14[7:7]<=0;end
else if(m14_7<1250)begin m14_7<=m14_7+1;end
else if(m14_7==1250)begin m14_7<=0;io14[7:7]<=~io14[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_8<=276;io14[8:8]<=1;end
else if(m14_8<1250)begin m14_8<=m14_8+1;end
else if(m14_8==1250)begin m14_8<=0;io14[8:8]<=~io14[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_9<=126;io14[9:9]<=0;end
else if(m14_9<1250)begin m14_9<=m14_9+1;end
else if(m14_9==1250)begin m14_9<=0;io14[9:9]<=~io14[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_10<=666;io14[10:10]<=0;end
else if(m14_10<1250)begin m14_10<=m14_10+1;end
else if(m14_10==1250)begin m14_10<=0;io14[10:10]<=~io14[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_11<=583;io14[11:11]<=1;end
else if(m14_11<1250)begin m14_11<=m14_11+1;end
else if(m14_11==1250)begin m14_11<=0;io14[11:11]<=~io14[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_12<=163;io14[12:12]<=0;end
else if(m14_12<1250)begin m14_12<=m14_12+1;end
else if(m14_12==1250)begin m14_12<=0;io14[12:12]<=~io14[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_13<=69;io14[13:13]<=0;end
else if(m14_13<1250)begin m14_13<=m14_13+1;end
else if(m14_13==1250)begin m14_13<=0;io14[13:13]<=~io14[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_14<=1069;io14[14:14]<=1;end
else if(m14_14<1250)begin m14_14<=m14_14+1;end
else if(m14_14==1250)begin m14_14<=0;io14[14:14]<=~io14[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_15<=35;io14[15:15]<=1;end
else if(m14_15<1250)begin m14_15<=m14_15+1;end
else if(m14_15==1250)begin m14_15<=0;io14[15:15]<=~io14[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_16<=185;io14[16:16]<=0;end
else if(m14_16<1250)begin m14_16<=m14_16+1;end
else if(m14_16==1250)begin m14_16<=0;io14[16:16]<=~io14[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_17<=662;io14[17:17]<=0;end
else if(m14_17<1250)begin m14_17<=m14_17+1;end
else if(m14_17==1250)begin m14_17<=0;io14[17:17]<=~io14[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_18<=767;io14[18:18]<=0;end
else if(m14_18<1250)begin m14_18<=m14_18+1;end
else if(m14_18==1250)begin m14_18<=0;io14[18:18]<=~io14[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_19<=490;io14[19:19]<=0;end
else if(m14_19<1250)begin m14_19<=m14_19+1;end
else if(m14_19==1250)begin m14_19<=0;io14[19:19]<=~io14[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_20<=256;io14[20:20]<=0;end
else if(m14_20<1250)begin m14_20<=m14_20+1;end
else if(m14_20==1250)begin m14_20<=0;io14[20:20]<=~io14[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_21<=283;io14[21:21]<=1;end
else if(m14_21<1250)begin m14_21<=m14_21+1;end
else if(m14_21==1250)begin m14_21<=0;io14[21:21]<=~io14[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_22<=828;io14[22:22]<=1;end
else if(m14_22<1250)begin m14_22<=m14_22+1;end
else if(m14_22==1250)begin m14_22<=0;io14[22:22]<=~io14[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_23<=762;io14[23:23]<=1;end
else if(m14_23<1250)begin m14_23<=m14_23+1;end
else if(m14_23==1250)begin m14_23<=0;io14[23:23]<=~io14[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m14_24<=729;io14[24:24]<=1;end
else if(m14_24<1250)begin m14_24<=m14_24+1;end
else if(m14_24==1250)begin m14_24<=0;io14[24:24]<=~io14[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_0<=145;io15[0:0]<=1;end
else if(m15_0<1250)begin m15_0<=m15_0+1;end
else if(m15_0==1250)begin m15_0<=0;io15[0:0]<=~io15[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_1<=398;io15[1:1]<=0;end
else if(m15_1<1250)begin m15_1<=m15_1+1;end
else if(m15_1==1250)begin m15_1<=0;io15[1:1]<=~io15[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_2<=309;io15[2:2]<=1;end
else if(m15_2<1250)begin m15_2<=m15_2+1;end
else if(m15_2==1250)begin m15_2<=0;io15[2:2]<=~io15[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_3<=860;io15[3:3]<=1;end
else if(m15_3<1250)begin m15_3<=m15_3+1;end
else if(m15_3==1250)begin m15_3<=0;io15[3:3]<=~io15[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_4<=756;io15[4:4]<=1;end
else if(m15_4<1250)begin m15_4<=m15_4+1;end
else if(m15_4==1250)begin m15_4<=0;io15[4:4]<=~io15[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_5<=46;io15[5:5]<=1;end
else if(m15_5<1250)begin m15_5<=m15_5+1;end
else if(m15_5==1250)begin m15_5<=0;io15[5:5]<=~io15[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_6<=1207;io15[6:6]<=0;end
else if(m15_6<1250)begin m15_6<=m15_6+1;end
else if(m15_6==1250)begin m15_6<=0;io15[6:6]<=~io15[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_7<=474;io15[7:7]<=0;end
else if(m15_7<1250)begin m15_7<=m15_7+1;end
else if(m15_7==1250)begin m15_7<=0;io15[7:7]<=~io15[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_8<=659;io15[8:8]<=1;end
else if(m15_8<1250)begin m15_8<=m15_8+1;end
else if(m15_8==1250)begin m15_8<=0;io15[8:8]<=~io15[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_9<=605;io15[9:9]<=0;end
else if(m15_9<1250)begin m15_9<=m15_9+1;end
else if(m15_9==1250)begin m15_9<=0;io15[9:9]<=~io15[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_10<=851;io15[10:10]<=0;end
else if(m15_10<1250)begin m15_10<=m15_10+1;end
else if(m15_10==1250)begin m15_10<=0;io15[10:10]<=~io15[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_11<=835;io15[11:11]<=1;end
else if(m15_11<1250)begin m15_11<=m15_11+1;end
else if(m15_11==1250)begin m15_11<=0;io15[11:11]<=~io15[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_12<=470;io15[12:12]<=0;end
else if(m15_12<1250)begin m15_12<=m15_12+1;end
else if(m15_12==1250)begin m15_12<=0;io15[12:12]<=~io15[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_13<=449;io15[13:13]<=0;end
else if(m15_13<1250)begin m15_13<=m15_13+1;end
else if(m15_13==1250)begin m15_13<=0;io15[13:13]<=~io15[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_14<=320;io15[14:14]<=0;end
else if(m15_14<1250)begin m15_14<=m15_14+1;end
else if(m15_14==1250)begin m15_14<=0;io15[14:14]<=~io15[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_15<=240;io15[15:15]<=1;end
else if(m15_15<1250)begin m15_15<=m15_15+1;end
else if(m15_15==1250)begin m15_15<=0;io15[15:15]<=~io15[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_16<=489;io15[16:16]<=0;end
else if(m15_16<1250)begin m15_16<=m15_16+1;end
else if(m15_16==1250)begin m15_16<=0;io15[16:16]<=~io15[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_17<=975;io15[17:17]<=0;end
else if(m15_17<1250)begin m15_17<=m15_17+1;end
else if(m15_17==1250)begin m15_17<=0;io15[17:17]<=~io15[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_18<=1156;io15[18:18]<=0;end
else if(m15_18<1250)begin m15_18<=m15_18+1;end
else if(m15_18==1250)begin m15_18<=0;io15[18:18]<=~io15[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_19<=924;io15[19:19]<=0;end
else if(m15_19<1250)begin m15_19<=m15_19+1;end
else if(m15_19==1250)begin m15_19<=0;io15[19:19]<=~io15[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_20<=485;io15[20:20]<=0;end
else if(m15_20<1250)begin m15_20<=m15_20+1;end
else if(m15_20==1250)begin m15_20<=0;io15[20:20]<=~io15[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_21<=453;io15[21:21]<=1;end
else if(m15_21<1250)begin m15_21<=m15_21+1;end
else if(m15_21==1250)begin m15_21<=0;io15[21:21]<=~io15[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_22<=1178;io15[22:22]<=1;end
else if(m15_22<1250)begin m15_22<=m15_22+1;end
else if(m15_22==1250)begin m15_22<=0;io15[22:22]<=~io15[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_23<=1137;io15[23:23]<=1;end
else if(m15_23<1250)begin m15_23<=m15_23+1;end
else if(m15_23==1250)begin m15_23<=0;io15[23:23]<=~io15[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m15_24<=1072;io15[24:24]<=1;end
else if(m15_24<1250)begin m15_24<=m15_24+1;end
else if(m15_24==1250)begin m15_24<=0;io15[24:24]<=~io15[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_0<=385;io16[0:0]<=1;end
else if(m16_0<1250)begin m16_0<=m16_0+1;end
else if(m16_0==1250)begin m16_0<=0;io16[0:0]<=~io16[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_1<=581;io16[1:1]<=0;end
else if(m16_1<1250)begin m16_1<=m16_1+1;end
else if(m16_1==1250)begin m16_1<=0;io16[1:1]<=~io16[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_2<=461;io16[2:2]<=1;end
else if(m16_2<1250)begin m16_2<=m16_2+1;end
else if(m16_2==1250)begin m16_2<=0;io16[2:2]<=~io16[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_3<=933;io16[3:3]<=1;end
else if(m16_3<1250)begin m16_3<=m16_3+1;end
else if(m16_3==1250)begin m16_3<=0;io16[3:3]<=~io16[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_4<=785;io16[4:4]<=1;end
else if(m16_4<1250)begin m16_4<=m16_4+1;end
else if(m16_4==1250)begin m16_4<=0;io16[4:4]<=~io16[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_5<=89;io16[5:5]<=1;end
else if(m16_5<1250)begin m16_5<=m16_5+1;end
else if(m16_5==1250)begin m16_5<=0;io16[5:5]<=~io16[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_6<=87;io16[6:6]<=1;end
else if(m16_6<1250)begin m16_6<=m16_6+1;end
else if(m16_6==1250)begin m16_6<=0;io16[6:6]<=~io16[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_7<=652;io16[7:7]<=0;end
else if(m16_7<1250)begin m16_7<=m16_7+1;end
else if(m16_7==1250)begin m16_7<=0;io16[7:7]<=~io16[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_8<=937;io16[8:8]<=1;end
else if(m16_8<1250)begin m16_8<=m16_8+1;end
else if(m16_8==1250)begin m16_8<=0;io16[8:8]<=~io16[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_9<=973;io16[9:9]<=0;end
else if(m16_9<1250)begin m16_9<=m16_9+1;end
else if(m16_9==1250)begin m16_9<=0;io16[9:9]<=~io16[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_10<=964;io16[10:10]<=0;end
else if(m16_10<1250)begin m16_10<=m16_10+1;end
else if(m16_10==1250)begin m16_10<=0;io16[10:10]<=~io16[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_11<=1015;io16[11:11]<=1;end
else if(m16_11<1250)begin m16_11<=m16_11+1;end
else if(m16_11==1250)begin m16_11<=0;io16[11:11]<=~io16[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_12<=721;io16[12:12]<=0;end
else if(m16_12<1250)begin m16_12<=m16_12+1;end
else if(m16_12==1250)begin m16_12<=0;io16[12:12]<=~io16[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_13<=778;io16[13:13]<=0;end
else if(m16_13<1250)begin m16_13<=m16_13+1;end
else if(m16_13==1250)begin m16_13<=0;io16[13:13]<=~io16[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_14<=741;io16[14:14]<=0;end
else if(m16_14<1250)begin m16_14<=m16_14+1;end
else if(m16_14==1250)begin m16_14<=0;io16[14:14]<=~io16[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_15<=408;io16[15:15]<=1;end
else if(m16_15<1250)begin m16_15<=m16_15+1;end
else if(m16_15==1250)begin m16_15<=0;io16[15:15]<=~io16[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_16<=754;io16[16:16]<=0;end
else if(m16_16<1250)begin m16_16<=m16_16+1;end
else if(m16_16==1250)begin m16_16<=0;io16[16:16]<=~io16[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_17<=36;io16[17:17]<=1;end
else if(m16_17<1250)begin m16_17<=m16_17+1;end
else if(m16_17==1250)begin m16_17<=0;io16[17:17]<=~io16[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_18<=308;io16[18:18]<=1;end
else if(m16_18<1250)begin m16_18<=m16_18+1;end
else if(m16_18==1250)begin m16_18<=0;io16[18:18]<=~io16[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_19<=29;io16[19:19]<=1;end
else if(m16_19<1250)begin m16_19<=m16_19+1;end
else if(m16_19==1250)begin m16_19<=0;io16[19:19]<=~io16[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_20<=768;io16[20:20]<=0;end
else if(m16_20<1250)begin m16_20<=m16_20+1;end
else if(m16_20==1250)begin m16_20<=0;io16[20:20]<=~io16[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_21<=650;io16[21:21]<=1;end
else if(m16_21<1250)begin m16_21<=m16_21+1;end
else if(m16_21==1250)begin m16_21<=0;io16[21:21]<=~io16[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_22<=359;io16[22:22]<=0;end
else if(m16_22<1250)begin m16_22<=m16_22+1;end
else if(m16_22==1250)begin m16_22<=0;io16[22:22]<=~io16[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_23<=329;io16[23:23]<=0;end
else if(m16_23<1250)begin m16_23<=m16_23+1;end
else if(m16_23==1250)begin m16_23<=0;io16[23:23]<=~io16[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m16_24<=176;io16[24:24]<=0;end
else if(m16_24<1250)begin m16_24<=m16_24+1;end
else if(m16_24==1250)begin m16_24<=0;io16[24:24]<=~io16[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_0<=385;io17[0:0]<=1;end
else if(m17_0<1250)begin m17_0<=m17_0+1;end
else if(m17_0==1250)begin m17_0<=0;io17[0:0]<=~io17[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_1<=581;io17[1:1]<=0;end
else if(m17_1<1250)begin m17_1<=m17_1+1;end
else if(m17_1==1250)begin m17_1<=0;io17[1:1]<=~io17[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_2<=461;io17[2:2]<=1;end
else if(m17_2<1250)begin m17_2<=m17_2+1;end
else if(m17_2==1250)begin m17_2<=0;io17[2:2]<=~io17[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_3<=933;io17[3:3]<=1;end
else if(m17_3<1250)begin m17_3<=m17_3+1;end
else if(m17_3==1250)begin m17_3<=0;io17[3:3]<=~io17[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_4<=785;io17[4:4]<=1;end
else if(m17_4<1250)begin m17_4<=m17_4+1;end
else if(m17_4==1250)begin m17_4<=0;io17[4:4]<=~io17[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_5<=89;io17[5:5]<=1;end
else if(m17_5<1250)begin m17_5<=m17_5+1;end
else if(m17_5==1250)begin m17_5<=0;io17[5:5]<=~io17[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_6<=87;io17[6:6]<=1;end
else if(m17_6<1250)begin m17_6<=m17_6+1;end
else if(m17_6==1250)begin m17_6<=0;io17[6:6]<=~io17[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_7<=652;io17[7:7]<=0;end
else if(m17_7<1250)begin m17_7<=m17_7+1;end
else if(m17_7==1250)begin m17_7<=0;io17[7:7]<=~io17[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_8<=937;io17[8:8]<=1;end
else if(m17_8<1250)begin m17_8<=m17_8+1;end
else if(m17_8==1250)begin m17_8<=0;io17[8:8]<=~io17[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_9<=973;io17[9:9]<=0;end
else if(m17_9<1250)begin m17_9<=m17_9+1;end
else if(m17_9==1250)begin m17_9<=0;io17[9:9]<=~io17[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_10<=964;io17[10:10]<=0;end
else if(m17_10<1250)begin m17_10<=m17_10+1;end
else if(m17_10==1250)begin m17_10<=0;io17[10:10]<=~io17[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_11<=1015;io17[11:11]<=1;end
else if(m17_11<1250)begin m17_11<=m17_11+1;end
else if(m17_11==1250)begin m17_11<=0;io17[11:11]<=~io17[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_12<=721;io17[12:12]<=0;end
else if(m17_12<1250)begin m17_12<=m17_12+1;end
else if(m17_12==1250)begin m17_12<=0;io17[12:12]<=~io17[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_13<=778;io17[13:13]<=0;end
else if(m17_13<1250)begin m17_13<=m17_13+1;end
else if(m17_13==1250)begin m17_13<=0;io17[13:13]<=~io17[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_14<=741;io17[14:14]<=0;end
else if(m17_14<1250)begin m17_14<=m17_14+1;end
else if(m17_14==1250)begin m17_14<=0;io17[14:14]<=~io17[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_15<=408;io17[15:15]<=1;end
else if(m17_15<1250)begin m17_15<=m17_15+1;end
else if(m17_15==1250)begin m17_15<=0;io17[15:15]<=~io17[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_16<=754;io17[16:16]<=0;end
else if(m17_16<1250)begin m17_16<=m17_16+1;end
else if(m17_16==1250)begin m17_16<=0;io17[16:16]<=~io17[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_17<=36;io17[17:17]<=1;end
else if(m17_17<1250)begin m17_17<=m17_17+1;end
else if(m17_17==1250)begin m17_17<=0;io17[17:17]<=~io17[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_18<=308;io17[18:18]<=1;end
else if(m17_18<1250)begin m17_18<=m17_18+1;end
else if(m17_18==1250)begin m17_18<=0;io17[18:18]<=~io17[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_19<=29;io17[19:19]<=1;end
else if(m17_19<1250)begin m17_19<=m17_19+1;end
else if(m17_19==1250)begin m17_19<=0;io17[19:19]<=~io17[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_20<=768;io17[20:20]<=0;end
else if(m17_20<1250)begin m17_20<=m17_20+1;end
else if(m17_20==1250)begin m17_20<=0;io17[20:20]<=~io17[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_21<=650;io17[21:21]<=1;end
else if(m17_21<1250)begin m17_21<=m17_21+1;end
else if(m17_21==1250)begin m17_21<=0;io17[21:21]<=~io17[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_22<=359;io17[22:22]<=0;end
else if(m17_22<1250)begin m17_22<=m17_22+1;end
else if(m17_22==1250)begin m17_22<=0;io17[22:22]<=~io17[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_23<=329;io17[23:23]<=0;end
else if(m17_23<1250)begin m17_23<=m17_23+1;end
else if(m17_23==1250)begin m17_23<=0;io17[23:23]<=~io17[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m17_24<=176;io17[24:24]<=0;end
else if(m17_24<1250)begin m17_24<=m17_24+1;end
else if(m17_24==1250)begin m17_24<=0;io17[24:24]<=~io17[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_0<=344;io18[0:0]<=1;end
else if(m18_0<1250)begin m18_0<=m18_0+1;end
else if(m18_0==1250)begin m18_0<=0;io18[0:0]<=~io18[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_1<=431;io18[1:1]<=0;end
else if(m18_1<1250)begin m18_1<=m18_1+1;end
else if(m18_1==1250)begin m18_1<=0;io18[1:1]<=~io18[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_2<=296;io18[2:2]<=1;end
else if(m18_2<1250)begin m18_2<=m18_2+1;end
else if(m18_2==1250)begin m18_2<=0;io18[2:2]<=~io18[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_3<=706;io18[3:3]<=1;end
else if(m18_3<1250)begin m18_3<=m18_3+1;end
else if(m18_3==1250)begin m18_3<=0;io18[3:3]<=~io18[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_4<=472;io18[4:4]<=1;end
else if(m18_4<1250)begin m18_4<=m18_4+1;end
else if(m18_4==1250)begin m18_4<=0;io18[4:4]<=~io18[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_5<=1041;io18[5:5]<=0;end
else if(m18_5<1250)begin m18_5<=m18_5+1;end
else if(m18_5==1250)begin m18_5<=0;io18[5:5]<=~io18[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_6<=1068;io18[6:6]<=0;end
else if(m18_6<1250)begin m18_6<=m18_6+1;end
else if(m18_6==1250)begin m18_6<=0;io18[6:6]<=~io18[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_7<=457;io18[7:7]<=0;end
else if(m18_7<1250)begin m18_7<=m18_7+1;end
else if(m18_7==1250)begin m18_7<=0;io18[7:7]<=~io18[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_8<=848;io18[8:8]<=1;end
else if(m18_8<1250)begin m18_8<=m18_8+1;end
else if(m18_8==1250)begin m18_8<=0;io18[8:8]<=~io18[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_9<=896;io18[9:9]<=0;end
else if(m18_9<1250)begin m18_9<=m18_9+1;end
else if(m18_9==1250)begin m18_9<=0;io18[9:9]<=~io18[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_10<=665;io18[10:10]<=0;end
else if(m18_10<1250)begin m18_10<=m18_10+1;end
else if(m18_10==1250)begin m18_10<=0;io18[10:10]<=~io18[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_11<=736;io18[11:11]<=1;end
else if(m18_11<1250)begin m18_11<=m18_11+1;end
else if(m18_11==1250)begin m18_11<=0;io18[11:11]<=~io18[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_12<=528;io18[12:12]<=0;end
else if(m18_12<1250)begin m18_12<=m18_12+1;end
else if(m18_12==1250)begin m18_12<=0;io18[12:12]<=~io18[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_13<=676;io18[13:13]<=0;end
else if(m18_13<1250)begin m18_13<=m18_13+1;end
else if(m18_13==1250)begin m18_13<=0;io18[13:13]<=~io18[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_14<=659;io18[14:14]<=0;end
else if(m18_14<1250)begin m18_14<=m18_14+1;end
else if(m18_14==1250)begin m18_14<=0;io18[14:14]<=~io18[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_15<=85;io18[15:15]<=1;end
else if(m18_15<1250)begin m18_15<=m18_15+1;end
else if(m18_15==1250)begin m18_15<=0;io18[15:15]<=~io18[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_16<=515;io18[16:16]<=0;end
else if(m18_16<1250)begin m18_16<=m18_16+1;end
else if(m18_16==1250)begin m18_16<=0;io18[16:16]<=~io18[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_17<=1110;io18[17:17]<=0;end
else if(m18_17<1250)begin m18_17<=m18_17+1;end
else if(m18_17==1250)begin m18_17<=0;io18[17:17]<=~io18[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_18<=171;io18[18:18]<=1;end
else if(m18_18<1250)begin m18_18<=m18_18+1;end
else if(m18_18==1250)begin m18_18<=0;io18[18:18]<=~io18[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_19<=1195;io18[19:19]<=0;end
else if(m18_19<1250)begin m18_19<=m18_19+1;end
else if(m18_19==1250)begin m18_19<=0;io18[19:19]<=~io18[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_20<=479;io18[20:20]<=0;end
else if(m18_20<1250)begin m18_20<=m18_20+1;end
else if(m18_20==1250)begin m18_20<=0;io18[20:20]<=~io18[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_21<=416;io18[21:21]<=1;end
else if(m18_21<1250)begin m18_21<=m18_21+1;end
else if(m18_21==1250)begin m18_21<=0;io18[21:21]<=~io18[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_22<=192;io18[22:22]<=0;end
else if(m18_22<1250)begin m18_22<=m18_22+1;end
else if(m18_22==1250)begin m18_22<=0;io18[22:22]<=~io18[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_23<=197;io18[23:23]<=0;end
else if(m18_23<1250)begin m18_23<=m18_23+1;end
else if(m18_23==1250)begin m18_23<=0;io18[23:23]<=~io18[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m18_24<=227;io18[24:24]<=0;end
else if(m18_24<1250)begin m18_24<=m18_24+1;end
else if(m18_24==1250)begin m18_24<=0;io18[24:24]<=~io18[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_0<=597;io19[0:0]<=1;end
else if(m19_0<1250)begin m19_0<=m19_0+1;end
else if(m19_0==1250)begin m19_0<=0;io19[0:0]<=~io19[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_1<=619;io19[1:1]<=0;end
else if(m19_1<1250)begin m19_1<=m19_1+1;end
else if(m19_1==1250)begin m19_1<=0;io19[1:1]<=~io19[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_2<=488;io19[2:2]<=1;end
else if(m19_2<1250)begin m19_2<=m19_2+1;end
else if(m19_2==1250)begin m19_2<=0;io19[2:2]<=~io19[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_3<=828;io19[3:3]<=1;end
else if(m19_3<1250)begin m19_3<=m19_3+1;end
else if(m19_3==1250)begin m19_3<=0;io19[3:3]<=~io19[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_4<=574;io19[4:4]<=1;end
else if(m19_4<1250)begin m19_4<=m19_4+1;end
else if(m19_4==1250)begin m19_4<=0;io19[4:4]<=~io19[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_5<=1135;io19[5:5]<=0;end
else if(m19_5<1250)begin m19_5<=m19_5+1;end
else if(m19_5==1250)begin m19_5<=0;io19[5:5]<=~io19[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_6<=1195;io19[6:6]<=0;end
else if(m19_6<1250)begin m19_6<=m19_6+1;end
else if(m19_6==1250)begin m19_6<=0;io19[6:6]<=~io19[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_7<=625;io19[7:7]<=0;end
else if(m19_7<1250)begin m19_7<=m19_7+1;end
else if(m19_7==1250)begin m19_7<=0;io19[7:7]<=~io19[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_8<=1044;io19[8:8]<=1;end
else if(m19_8<1250)begin m19_8<=m19_8+1;end
else if(m19_8==1250)begin m19_8<=0;io19[8:8]<=~io19[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_9<=1094;io19[9:9]<=0;end
else if(m19_9<1250)begin m19_9<=m19_9+1;end
else if(m19_9==1250)begin m19_9<=0;io19[9:9]<=~io19[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_10<=757;io19[10:10]<=0;end
else if(m19_10<1250)begin m19_10<=m19_10+1;end
else if(m19_10==1250)begin m19_10<=0;io19[10:10]<=~io19[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_11<=870;io19[11:11]<=1;end
else if(m19_11<1250)begin m19_11<=m19_11+1;end
else if(m19_11==1250)begin m19_11<=0;io19[11:11]<=~io19[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_12<=700;io19[12:12]<=0;end
else if(m19_12<1250)begin m19_12<=m19_12+1;end
else if(m19_12==1250)begin m19_12<=0;io19[12:12]<=~io19[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_13<=870;io19[13:13]<=0;end
else if(m19_13<1250)begin m19_13<=m19_13+1;end
else if(m19_13==1250)begin m19_13<=0;io19[13:13]<=~io19[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_14<=830;io19[14:14]<=0;end
else if(m19_14<1250)begin m19_14<=m19_14+1;end
else if(m19_14==1250)begin m19_14<=0;io19[14:14]<=~io19[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_15<=175;io19[15:15]<=1;end
else if(m19_15<1250)begin m19_15<=m19_15+1;end
else if(m19_15==1250)begin m19_15<=0;io19[15:15]<=~io19[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_16<=635;io19[16:16]<=0;end
else if(m19_16<1250)begin m19_16<=m19_16+1;end
else if(m19_16==1250)begin m19_16<=0;io19[16:16]<=~io19[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_17<=49;io19[17:17]<=1;end
else if(m19_17<1250)begin m19_17<=m19_17+1;end
else if(m19_17==1250)begin m19_17<=0;io19[17:17]<=~io19[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_18<=357;io19[18:18]<=1;end
else if(m19_18<1250)begin m19_18<=m19_18+1;end
else if(m19_18==1250)begin m19_18<=0;io19[18:18]<=~io19[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_19<=186;io19[19:19]<=1;end
else if(m19_19<1250)begin m19_19<=m19_19+1;end
else if(m19_19==1250)begin m19_19<=0;io19[19:19]<=~io19[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_20<=591;io19[20:20]<=0;end
else if(m19_20<1250)begin m19_20<=m19_20+1;end
else if(m19_20==1250)begin m19_20<=0;io19[20:20]<=~io19[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_21<=580;io19[21:21]<=1;end
else if(m19_21<1250)begin m19_21<=m19_21+1;end
else if(m19_21==1250)begin m19_21<=0;io19[21:21]<=~io19[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_22<=358;io19[22:22]<=0;end
else if(m19_22<1250)begin m19_22<=m19_22+1;end
else if(m19_22==1250)begin m19_22<=0;io19[22:22]<=~io19[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_23<=406;io19[23:23]<=0;end
else if(m19_23<1250)begin m19_23<=m19_23+1;end
else if(m19_23==1250)begin m19_23<=0;io19[23:23]<=~io19[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m19_24<=485;io19[24:24]<=0;end
else if(m19_24<1250)begin m19_24<=m19_24+1;end
else if(m19_24==1250)begin m19_24<=0;io19[24:24]<=~io19[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_0<=1007;io20[0:0]<=0;end
else if(m20_0<1250)begin m20_0<=m20_0+1;end
else if(m20_0==1250)begin m20_0<=0;io20[0:0]<=~io20[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_1<=880;io20[1:1]<=1;end
else if(m20_1<1250)begin m20_1<=m20_1+1;end
else if(m20_1==1250)begin m20_1<=0;io20[1:1]<=~io20[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_2<=894;io20[2:2]<=0;end
else if(m20_2<1250)begin m20_2<=m20_2+1;end
else if(m20_2==1250)begin m20_2<=0;io20[2:2]<=~io20[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_3<=866;io20[3:3]<=1;end
else if(m20_3<1250)begin m20_3<=m20_3+1;end
else if(m20_3==1250)begin m20_3<=0;io20[3:3]<=~io20[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_4<=966;io20[4:4]<=0;end
else if(m20_4<1250)begin m20_4<=m20_4+1;end
else if(m20_4==1250)begin m20_4<=0;io20[4:4]<=~io20[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_5<=289;io20[5:5]<=0;end
else if(m20_5<1250)begin m20_5<=m20_5+1;end
else if(m20_5==1250)begin m20_5<=0;io20[5:5]<=~io20[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_6<=91;io20[6:6]<=1;end
else if(m20_6<1250)begin m20_6<=m20_6+1;end
else if(m20_6==1250)begin m20_6<=0;io20[6:6]<=~io20[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_7<=1041;io20[7:7]<=1;end
else if(m20_7<1250)begin m20_7<=m20_7+1;end
else if(m20_7==1250)begin m20_7<=0;io20[7:7]<=~io20[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_8<=98;io20[8:8]<=1;end
else if(m20_8<1250)begin m20_8<=m20_8+1;end
else if(m20_8==1250)begin m20_8<=0;io20[8:8]<=~io20[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_9<=289;io20[9:9]<=0;end
else if(m20_9<1250)begin m20_9<=m20_9+1;end
else if(m20_9==1250)begin m20_9<=0;io20[9:9]<=~io20[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_10<=1201;io20[10:10]<=1;end
else if(m20_10<1250)begin m20_10<=m20_10+1;end
else if(m20_10==1250)begin m20_10<=0;io20[10:10]<=~io20[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_11<=1185;io20[11:11]<=1;end
else if(m20_11<1250)begin m20_11<=m20_11+1;end
else if(m20_11==1250)begin m20_11<=0;io20[11:11]<=~io20[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_12<=1109;io20[12:12]<=1;end
else if(m20_12<1250)begin m20_12<=m20_12+1;end
else if(m20_12==1250)begin m20_12<=0;io20[12:12]<=~io20[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_13<=46;io20[13:13]<=0;end
else if(m20_13<1250)begin m20_13<=m20_13+1;end
else if(m20_13==1250)begin m20_13<=0;io20[13:13]<=~io20[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_14<=1229;io20[14:14]<=1;end
else if(m20_14<1250)begin m20_14<=m20_14+1;end
else if(m20_14==1250)begin m20_14<=0;io20[14:14]<=~io20[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_15<=570;io20[15:15]<=0;end
else if(m20_15<1250)begin m20_15<=m20_15+1;end
else if(m20_15==1250)begin m20_15<=0;io20[15:15]<=~io20[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_16<=702;io20[16:16]<=0;end
else if(m20_16<1250)begin m20_16<=m20_16+1;end
else if(m20_16==1250)begin m20_16<=0;io20[16:16]<=~io20[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_17<=459;io20[17:17]<=0;end
else if(m20_17<1250)begin m20_17<=m20_17+1;end
else if(m20_17==1250)begin m20_17<=0;io20[17:17]<=~io20[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_18<=605;io20[18:18]<=0;end
else if(m20_18<1250)begin m20_18<=m20_18+1;end
else if(m20_18==1250)begin m20_18<=0;io20[18:18]<=~io20[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_19<=633;io20[19:19]<=0;end
else if(m20_19<1250)begin m20_19<=m20_19+1;end
else if(m20_19==1250)begin m20_19<=0;io20[19:19]<=~io20[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_20<=962;io20[20:20]<=1;end
else if(m20_20<1250)begin m20_20<=m20_20+1;end
else if(m20_20==1250)begin m20_20<=0;io20[20:20]<=~io20[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_21<=904;io20[21:21]<=1;end
else if(m20_21<1250)begin m20_21<=m20_21+1;end
else if(m20_21==1250)begin m20_21<=0;io20[21:21]<=~io20[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_22<=768;io20[22:22]<=1;end
else if(m20_22<1250)begin m20_22<=m20_22+1;end
else if(m20_22==1250)begin m20_22<=0;io20[22:22]<=~io20[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_23<=800;io20[23:23]<=1;end
else if(m20_23<1250)begin m20_23<=m20_23+1;end
else if(m20_23==1250)begin m20_23<=0;io20[23:23]<=~io20[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m20_24<=914;io20[24:24]<=1;end
else if(m20_24<1250)begin m20_24<=m20_24+1;end
else if(m20_24==1250)begin m20_24<=0;io20[24:24]<=~io20[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_0<=513;io21[0:0]<=1;end
else if(m21_0<1250)begin m21_0<=m21_0+1;end
else if(m21_0==1250)begin m21_0<=0;io21[0:0]<=~io21[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_1<=720;io21[1:1]<=1;end
else if(m21_1<1250)begin m21_1<=m21_1+1;end
else if(m21_1==1250)begin m21_1<=0;io21[1:1]<=~io21[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_2<=296;io21[2:2]<=1;end
else if(m21_2<1250)begin m21_2<=m21_2+1;end
else if(m21_2==1250)begin m21_2<=0;io21[2:2]<=~io21[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_3<=417;io21[3:3]<=0;end
else if(m21_3<1250)begin m21_3<=m21_3+1;end
else if(m21_3==1250)begin m21_3<=0;io21[3:3]<=~io21[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_4<=302;io21[4:4]<=1;end
else if(m21_4<1250)begin m21_4<=m21_4+1;end
else if(m21_4==1250)begin m21_4<=0;io21[4:4]<=~io21[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_5<=896;io21[5:5]<=0;end
else if(m21_5<1250)begin m21_5<=m21_5+1;end
else if(m21_5==1250)begin m21_5<=0;io21[5:5]<=~io21[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_6<=841;io21[6:6]<=1;end
else if(m21_6<1250)begin m21_6<=m21_6+1;end
else if(m21_6==1250)begin m21_6<=0;io21[6:6]<=~io21[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_7<=457;io21[7:7]<=0;end
else if(m21_7<1250)begin m21_7<=m21_7+1;end
else if(m21_7==1250)begin m21_7<=0;io21[7:7]<=~io21[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_8<=1075;io21[8:8]<=0;end
else if(m21_8<1250)begin m21_8<=m21_8+1;end
else if(m21_8==1250)begin m21_8<=0;io21[8:8]<=~io21[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_9<=1041;io21[9:9]<=0;end
else if(m21_9<1250)begin m21_9<=m21_9+1;end
else if(m21_9==1250)begin m21_9<=0;io21[9:9]<=~io21[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_10<=632;io21[10:10]<=0;end
else if(m21_10<1250)begin m21_10<=m21_10+1;end
else if(m21_10==1250)begin m21_10<=0;io21[10:10]<=~io21[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_11<=565;io21[11:11]<=0;end
else if(m21_11<1250)begin m21_11<=m21_11+1;end
else if(m21_11==1250)begin m21_11<=0;io21[11:11]<=~io21[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_12<=528;io21[12:12]<=0;end
else if(m21_12<1250)begin m21_12<=m21_12+1;end
else if(m21_12==1250)begin m21_12<=0;io21[12:12]<=~io21[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_13<=848;io21[13:13]<=1;end
else if(m21_13<1250)begin m21_13<=m21_13+1;end
else if(m21_13==1250)begin m21_13<=0;io21[13:13]<=~io21[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_14<=693;io21[14:14]<=0;end
else if(m21_14<1250)begin m21_14<=m21_14+1;end
else if(m21_14==1250)begin m21_14<=0;io21[14:14]<=~io21[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_15<=1132;io21[15:15]<=0;end
else if(m21_15<1250)begin m21_15<=m21_15+1;end
else if(m21_15==1250)begin m21_15<=0;io21[15:15]<=~io21[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_16<=268;io21[16:16]<=1;end
else if(m21_16<1250)begin m21_16<=m21_16+1;end
else if(m21_16==1250)begin m21_16<=0;io21[16:16]<=~io21[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_17<=1110;io21[17:17]<=0;end
else if(m21_17<1250)begin m21_17<=m21_17+1;end
else if(m21_17==1250)begin m21_17<=0;io21[17:17]<=~io21[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_18<=418;io21[18:18]<=0;end
else if(m21_18<1250)begin m21_18<=m21_18+1;end
else if(m21_18==1250)begin m21_18<=0;io21[18:18]<=~io21[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_19<=147;io21[19:19]<=1;end
else if(m21_19<1250)begin m21_19<=m21_19+1;end
else if(m21_19==1250)begin m21_19<=0;io21[19:19]<=~io21[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_20<=275;io21[20:20]<=0;end
else if(m21_20<1250)begin m21_20<=m21_20+1;end
else if(m21_20==1250)begin m21_20<=0;io21[20:20]<=~io21[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_21<=301;io21[21:21]<=0;end
else if(m21_21<1250)begin m21_21<=m21_21+1;end
else if(m21_21==1250)begin m21_21<=0;io21[21:21]<=~io21[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_22<=192;io21[22:22]<=0;end
else if(m21_22<1250)begin m21_22<=m21_22+1;end
else if(m21_22==1250)begin m21_22<=0;io21[22:22]<=~io21[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_23<=311;io21[23:23]<=1;end
else if(m21_23<1250)begin m21_23<=m21_23+1;end
else if(m21_23==1250)begin m21_23<=0;io21[23:23]<=~io21[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m21_24<=431;io21[24:24]<=0;end
else if(m21_24<1250)begin m21_24<=m21_24+1;end
else if(m21_24==1250)begin m21_24<=0;io21[24:24]<=~io21[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_0<=513;io22[0:0]<=1;end
else if(m22_0<1250)begin m22_0<=m22_0+1;end
else if(m22_0==1250)begin m22_0<=0;io22[0:0]<=~io22[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_1<=720;io22[1:1]<=1;end
else if(m22_1<1250)begin m22_1<=m22_1+1;end
else if(m22_1==1250)begin m22_1<=0;io22[1:1]<=~io22[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_2<=296;io22[2:2]<=1;end
else if(m22_2<1250)begin m22_2<=m22_2+1;end
else if(m22_2==1250)begin m22_2<=0;io22[2:2]<=~io22[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_3<=417;io22[3:3]<=0;end
else if(m22_3<1250)begin m22_3<=m22_3+1;end
else if(m22_3==1250)begin m22_3<=0;io22[3:3]<=~io22[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_4<=302;io22[4:4]<=1;end
else if(m22_4<1250)begin m22_4<=m22_4+1;end
else if(m22_4==1250)begin m22_4<=0;io22[4:4]<=~io22[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_5<=896;io22[5:5]<=0;end
else if(m22_5<1250)begin m22_5<=m22_5+1;end
else if(m22_5==1250)begin m22_5<=0;io22[5:5]<=~io22[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_6<=841;io22[6:6]<=1;end
else if(m22_6<1250)begin m22_6<=m22_6+1;end
else if(m22_6==1250)begin m22_6<=0;io22[6:6]<=~io22[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_7<=457;io22[7:7]<=0;end
else if(m22_7<1250)begin m22_7<=m22_7+1;end
else if(m22_7==1250)begin m22_7<=0;io22[7:7]<=~io22[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_8<=1075;io22[8:8]<=0;end
else if(m22_8<1250)begin m22_8<=m22_8+1;end
else if(m22_8==1250)begin m22_8<=0;io22[8:8]<=~io22[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_9<=1041;io22[9:9]<=0;end
else if(m22_9<1250)begin m22_9<=m22_9+1;end
else if(m22_9==1250)begin m22_9<=0;io22[9:9]<=~io22[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_10<=632;io22[10:10]<=0;end
else if(m22_10<1250)begin m22_10<=m22_10+1;end
else if(m22_10==1250)begin m22_10<=0;io22[10:10]<=~io22[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_11<=565;io22[11:11]<=0;end
else if(m22_11<1250)begin m22_11<=m22_11+1;end
else if(m22_11==1250)begin m22_11<=0;io22[11:11]<=~io22[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_12<=528;io22[12:12]<=0;end
else if(m22_12<1250)begin m22_12<=m22_12+1;end
else if(m22_12==1250)begin m22_12<=0;io22[12:12]<=~io22[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_13<=848;io22[13:13]<=1;end
else if(m22_13<1250)begin m22_13<=m22_13+1;end
else if(m22_13==1250)begin m22_13<=0;io22[13:13]<=~io22[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_14<=693;io22[14:14]<=0;end
else if(m22_14<1250)begin m22_14<=m22_14+1;end
else if(m22_14==1250)begin m22_14<=0;io22[14:14]<=~io22[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_15<=1132;io22[15:15]<=0;end
else if(m22_15<1250)begin m22_15<=m22_15+1;end
else if(m22_15==1250)begin m22_15<=0;io22[15:15]<=~io22[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_16<=268;io22[16:16]<=1;end
else if(m22_16<1250)begin m22_16<=m22_16+1;end
else if(m22_16==1250)begin m22_16<=0;io22[16:16]<=~io22[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_17<=1110;io22[17:17]<=0;end
else if(m22_17<1250)begin m22_17<=m22_17+1;end
else if(m22_17==1250)begin m22_17<=0;io22[17:17]<=~io22[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_18<=418;io22[18:18]<=0;end
else if(m22_18<1250)begin m22_18<=m22_18+1;end
else if(m22_18==1250)begin m22_18<=0;io22[18:18]<=~io22[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_19<=147;io22[19:19]<=1;end
else if(m22_19<1250)begin m22_19<=m22_19+1;end
else if(m22_19==1250)begin m22_19<=0;io22[19:19]<=~io22[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_20<=275;io22[20:20]<=0;end
else if(m22_20<1250)begin m22_20<=m22_20+1;end
else if(m22_20==1250)begin m22_20<=0;io22[20:20]<=~io22[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_21<=301;io22[21:21]<=0;end
else if(m22_21<1250)begin m22_21<=m22_21+1;end
else if(m22_21==1250)begin m22_21<=0;io22[21:21]<=~io22[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_22<=192;io22[22:22]<=0;end
else if(m22_22<1250)begin m22_22<=m22_22+1;end
else if(m22_22==1250)begin m22_22<=0;io22[22:22]<=~io22[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_23<=311;io22[23:23]<=1;end
else if(m22_23<1250)begin m22_23<=m22_23+1;end
else if(m22_23==1250)begin m22_23<=0;io22[23:23]<=~io22[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m22_24<=431;io22[24:24]<=0;end
else if(m22_24<1250)begin m22_24<=m22_24+1;end
else if(m22_24==1250)begin m22_24<=0;io22[24:24]<=~io22[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_0<=629;io23[0:0]<=1;end
else if(m23_0<1250)begin m23_0<=m23_0+1;end
else if(m23_0==1250)begin m23_0<=0;io23[0:0]<=~io23[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_1<=771;io23[1:1]<=1;end
else if(m23_1<1250)begin m23_1<=m23_1+1;end
else if(m23_1==1250)begin m23_1<=0;io23[1:1]<=~io23[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_2<=253;io23[2:2]<=1;end
else if(m23_2<1250)begin m23_2<=m23_2+1;end
else if(m23_2==1250)begin m23_2<=0;io23[2:2]<=~io23[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_3<=350;io23[3:3]<=0;end
else if(m23_3<1250)begin m23_3<=m23_3+1;end
else if(m23_3==1250)begin m23_3<=0;io23[3:3]<=~io23[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_4<=113;io23[4:4]<=1;end
else if(m23_4<1250)begin m23_4<=m23_4+1;end
else if(m23_4==1250)begin m23_4<=0;io23[4:4]<=~io23[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_5<=668;io23[5:5]<=0;end
else if(m23_5<1250)begin m23_5<=m23_5+1;end
else if(m23_5==1250)begin m23_5<=0;io23[5:5]<=~io23[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_6<=671;io23[6:6]<=1;end
else if(m23_6<1250)begin m23_6<=m23_6+1;end
else if(m23_6==1250)begin m23_6<=0;io23[6:6]<=~io23[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_7<=376;io23[7:7]<=0;end
else if(m23_7<1250)begin m23_7<=m23_7+1;end
else if(m23_7==1250)begin m23_7<=0;io23[7:7]<=~io23[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_8<=1074;io23[8:8]<=0;end
else if(m23_8<1250)begin m23_8<=m23_8+1;end
else if(m23_8==1250)begin m23_8<=0;io23[8:8]<=~io23[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_9<=1087;io23[9:9]<=0;end
else if(m23_9<1250)begin m23_9<=m23_9+1;end
else if(m23_9==1250)begin m23_9<=0;io23[9:9]<=~io23[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_10<=354;io23[10:10]<=0;end
else if(m23_10<1250)begin m23_10<=m23_10+1;end
else if(m23_10==1250)begin m23_10<=0;io23[10:10]<=~io23[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_11<=340;io23[11:11]<=0;end
else if(m23_11<1250)begin m23_11<=m23_11+1;end
else if(m23_11==1250)begin m23_11<=0;io23[11:11]<=~io23[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_12<=383;io23[12:12]<=0;end
else if(m23_12<1250)begin m23_12<=m23_12+1;end
else if(m23_12==1250)begin m23_12<=0;io23[12:12]<=~io23[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_13<=790;io23[13:13]<=1;end
else if(m23_13<1250)begin m23_13<=m23_13+1;end
else if(m23_13==1250)begin m23_13<=0;io23[13:13]<=~io23[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_14<=669;io23[14:14]<=0;end
else if(m23_14<1250)begin m23_14<=m23_14+1;end
else if(m23_14==1250)begin m23_14<=0;io23[14:14]<=~io23[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_15<=872;io23[15:15]<=0;end
else if(m23_15<1250)begin m23_15<=m23_15+1;end
else if(m23_15==1250)begin m23_15<=0;io23[15:15]<=~io23[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_16<=1244;io23[16:16]<=0;end
else if(m23_16<1250)begin m23_16<=m23_16+1;end
else if(m23_16==1250)begin m23_16<=0;io23[16:16]<=~io23[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_17<=895;io23[17:17]<=0;end
else if(m23_17<1250)begin m23_17<=m23_17+1;end
else if(m23_17==1250)begin m23_17<=0;io23[17:17]<=~io23[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_18<=290;io23[18:18]<=0;end
else if(m23_18<1250)begin m23_18<=m23_18+1;end
else if(m23_18==1250)begin m23_18<=0;io23[18:18]<=~io23[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_19<=92;io23[19:19]<=1;end
else if(m23_19<1250)begin m23_19<=m23_19+1;end
else if(m23_19==1250)begin m23_19<=0;io23[19:19]<=~io23[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_20<=1122;io23[20:20]<=1;end
else if(m23_20<1250)begin m23_20<=m23_20+1;end
else if(m23_20==1250)begin m23_20<=0;io23[20:20]<=~io23[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_21<=1212;io23[21:21]<=1;end
else if(m23_21<1250)begin m23_21<=m23_21+1;end
else if(m23_21==1250)begin m23_21<=0;io23[21:21]<=~io23[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_22<=1143;io23[22:22]<=1;end
else if(m23_22<1250)begin m23_22<=m23_22+1;end
else if(m23_22==1250)begin m23_22<=0;io23[22:22]<=~io23[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_23<=183;io23[23:23]<=1;end
else if(m23_23<1250)begin m23_23<=m23_23+1;end
else if(m23_23==1250)begin m23_23<=0;io23[23:23]<=~io23[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m23_24<=273;io23[24:24]<=0;end
else if(m23_24<1250)begin m23_24<=m23_24+1;end
else if(m23_24==1250)begin m23_24<=0;io23[24:24]<=~io23[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_0<=798;io24[0:0]<=1;end
else if(m24_0<1250)begin m24_0<=m24_0+1;end
else if(m24_0==1250)begin m24_0<=0;io24[0:0]<=~io24[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_1<=874;io24[1:1]<=1;end
else if(m24_1<1250)begin m24_1<=m24_1+1;end
else if(m24_1==1250)begin m24_1<=0;io24[1:1]<=~io24[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_2<=309;io24[2:2]<=1;end
else if(m24_2<1250)begin m24_2<=m24_2+1;end
else if(m24_2==1250)begin m24_2<=0;io24[2:2]<=~io24[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_3<=384;io24[3:3]<=0;end
else if(m24_3<1250)begin m24_3<=m24_3+1;end
else if(m24_3==1250)begin m24_3<=0;io24[3:3]<=~io24[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_4<=103;io24[4:4]<=1;end
else if(m24_4<1250)begin m24_4<=m24_4+1;end
else if(m24_4==1250)begin m24_4<=0;io24[4:4]<=~io24[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_5<=605;io24[5:5]<=0;end
else if(m24_5<1250)begin m24_5<=m24_5+1;end
else if(m24_5==1250)begin m24_5<=0;io24[5:5]<=~io24[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_6<=652;io24[6:6]<=1;end
else if(m24_6<1250)begin m24_6<=m24_6+1;end
else if(m24_6==1250)begin m24_6<=0;io24[6:6]<=~io24[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_7<=474;io24[7:7]<=0;end
else if(m24_7<1250)begin m24_7<=m24_7+1;end
else if(m24_7==1250)begin m24_7<=0;io24[7:7]<=~io24[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_8<=1214;io24[8:8]<=0;end
else if(m24_8<1250)begin m24_8<=m24_8+1;end
else if(m24_8==1250)begin m24_8<=0;io24[8:8]<=~io24[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_9<=46;io24[9:9]<=1;end
else if(m24_9<1250)begin m24_9<=m24_9+1;end
else if(m24_9==1250)begin m24_9<=0;io24[9:9]<=~io24[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_10<=292;io24[10:10]<=0;end
else if(m24_10<1250)begin m24_10<=m24_10+1;end
else if(m24_10==1250)begin m24_10<=0;io24[10:10]<=~io24[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_11<=338;io24[11:11]<=0;end
else if(m24_11<1250)begin m24_11<=m24_11+1;end
else if(m24_11==1250)begin m24_11<=0;io24[11:11]<=~io24[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_12<=470;io24[12:12]<=0;end
else if(m24_12<1250)begin m24_12<=m24_12+1;end
else if(m24_12==1250)begin m24_12<=0;io24[12:12]<=~io24[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_13<=946;io24[13:13]<=1;end
else if(m24_13<1250)begin m24_13<=m24_13+1;end
else if(m24_13==1250)begin m24_13<=0;io24[13:13]<=~io24[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_14<=879;io24[14:14]<=0;end
else if(m24_14<1250)begin m24_14<=m24_14+1;end
else if(m24_14==1250)begin m24_14<=0;io24[14:14]<=~io24[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_15<=862;io24[15:15]<=0;end
else if(m24_15<1250)begin m24_15<=m24_15+1;end
else if(m24_15==1250)begin m24_15<=0;io24[15:15]<=~io24[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_16<=3;io24[16:16]<=1;end
else if(m24_16<1250)begin m24_16<=m24_16+1;end
else if(m24_16==1250)begin m24_16<=0;io24[16:16]<=~io24[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_17<=975;io24[17:17]<=0;end
else if(m24_17<1250)begin m24_17<=m24_17+1;end
else if(m24_17==1250)begin m24_17<=0;io24[17:17]<=~io24[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_18<=392;io24[18:18]<=0;end
else if(m24_18<1250)begin m24_18<=m24_18+1;end
else if(m24_18==1250)begin m24_18<=0;io24[18:18]<=~io24[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_19<=302;io24[19:19]<=1;end
else if(m24_19<1250)begin m24_19<=m24_19+1;end
else if(m24_19==1250)begin m24_19<=0;io24[19:19]<=~io24[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_20<=1120;io24[20:20]<=1;end
else if(m24_20<1250)begin m24_20<=m24_20+1;end
else if(m24_20==1250)begin m24_20<=0;io24[20:20]<=~io24[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_21<=1241;io24[21:21]<=1;end
else if(m24_21<1250)begin m24_21<=m24_21+1;end
else if(m24_21==1250)begin m24_21<=0;io24[21:21]<=~io24[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_22<=1178;io24[22:22]<=1;end
else if(m24_22<1250)begin m24_22<=m24_22+1;end
else if(m24_22==1250)begin m24_22<=0;io24[22:22]<=~io24[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_23<=349;io24[23:23]<=1;end
else if(m24_23<1250)begin m24_23<=m24_23+1;end
else if(m24_23==1250)begin m24_23<=0;io24[23:23]<=~io24[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m24_24<=436;io24[24:24]<=0;end
else if(m24_24<1250)begin m24_24<=m24_24+1;end
else if(m24_24==1250)begin m24_24<=0;io24[24:24]<=~io24[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_0<=896;io25[0:0]<=1;end
else if(m25_0<1250)begin m25_0<=m25_0+1;end
else if(m25_0==1250)begin m25_0<=0;io25[0:0]<=~io25[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_1<=1001;io25[1:1]<=1;end
else if(m25_1<1250)begin m25_1<=m25_1+1;end
else if(m25_1==1250)begin m25_1<=0;io25[1:1]<=~io25[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_2<=407;io25[2:2]<=1;end
else if(m25_2<1250)begin m25_2<=m25_2+1;end
else if(m25_2==1250)begin m25_2<=0;io25[2:2]<=~io25[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_3<=493;io25[3:3]<=0;end
else if(m25_3<1250)begin m25_3<=m25_3+1;end
else if(m25_3==1250)begin m25_3<=0;io25[3:3]<=~io25[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_4<=164;io25[4:4]<=1;end
else if(m25_4<1250)begin m25_4<=m25_4+1;end
else if(m25_4==1250)begin m25_4<=0;io25[4:4]<=~io25[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_5<=648;io25[5:5]<=0;end
else if(m25_5<1250)begin m25_5<=m25_5+1;end
else if(m25_5==1250)begin m25_5<=0;io25[5:5]<=~io25[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_6<=719;io25[6:6]<=1;end
else if(m25_6<1250)begin m25_6<=m25_6+1;end
else if(m25_6==1250)begin m25_6<=0;io25[6:6]<=~io25[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_7<=534;io25[7:7]<=0;end
else if(m25_7<1250)begin m25_7<=m25_7+1;end
else if(m25_7==1250)begin m25_7<=0;io25[7:7]<=~io25[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_8<=1248;io25[8:8]<=0;end
else if(m25_8<1250)begin m25_8<=m25_8+1;end
else if(m25_8==1250)begin m25_8<=0;io25[8:8]<=~io25[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_9<=119;io25[9:9]<=1;end
else if(m25_9<1250)begin m25_9<=m25_9+1;end
else if(m25_9==1250)begin m25_9<=0;io25[9:9]<=~io25[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_10<=223;io25[10:10]<=0;end
else if(m25_10<1250)begin m25_10<=m25_10+1;end
else if(m25_10==1250)begin m25_10<=0;io25[10:10]<=~io25[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_11<=310;io25[11:11]<=0;end
else if(m25_11<1250)begin m25_11<=m25_11+1;end
else if(m25_11==1250)begin m25_11<=0;io25[11:11]<=~io25[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_12<=428;io25[12:12]<=0;end
else if(m25_12<1250)begin m25_12<=m25_12+1;end
else if(m25_12==1250)begin m25_12<=0;io25[12:12]<=~io25[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_13<=923;io25[13:13]<=1;end
else if(m25_13<1250)begin m25_13<=m25_13+1;end
else if(m25_13==1250)begin m25_13<=0;io25[13:13]<=~io25[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_14<=871;io25[14:14]<=0;end
else if(m25_14<1250)begin m25_14<=m25_14+1;end
else if(m25_14==1250)begin m25_14<=0;io25[14:14]<=~io25[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_15<=828;io25[15:15]<=0;end
else if(m25_15<1250)begin m25_15<=m25_15+1;end
else if(m25_15==1250)begin m25_15<=0;io25[15:15]<=~io25[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_16<=1154;io25[16:16]<=0;end
else if(m25_16<1250)begin m25_16<=m25_16+1;end
else if(m25_16==1250)begin m25_16<=0;io25[16:16]<=~io25[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_17<=910;io25[17:17]<=0;end
else if(m25_17<1250)begin m25_17<=m25_17+1;end
else if(m25_17==1250)begin m25_17<=0;io25[17:17]<=~io25[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_18<=336;io25[18:18]<=0;end
else if(m25_18<1250)begin m25_18<=m25_18+1;end
else if(m25_18==1250)begin m25_18<=0;io25[18:18]<=~io25[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_19<=237;io25[19:19]<=1;end
else if(m25_19<1250)begin m25_19<=m25_19+1;end
else if(m25_19==1250)begin m25_19<=0;io25[19:19]<=~io25[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_20<=1032;io25[20:20]<=1;end
else if(m25_20<1250)begin m25_20<=m25_20+1;end
else if(m25_20==1250)begin m25_20<=0;io25[20:20]<=~io25[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_21<=1112;io25[21:21]<=1;end
else if(m25_21<1250)begin m25_21<=m25_21+1;end
else if(m25_21==1250)begin m25_21<=0;io25[21:21]<=~io25[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_22<=1045;io25[22:22]<=1;end
else if(m25_22<1250)begin m25_22<=m25_22+1;end
else if(m25_22==1250)begin m25_22<=0;io25[22:22]<=~io25[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_23<=263;io25[23:23]<=1;end
else if(m25_23<1250)begin m25_23<=m25_23+1;end
else if(m25_23==1250)begin m25_23<=0;io25[23:23]<=~io25[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m25_24<=309;io25[24:24]<=0;end
else if(m25_24<1250)begin m25_24<=m25_24+1;end
else if(m25_24==1250)begin m25_24<=0;io25[24:24]<=~io25[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_0<=896;io26[0:0]<=1;end
else if(m26_0<1250)begin m26_0<=m26_0+1;end
else if(m26_0==1250)begin m26_0<=0;io26[0:0]<=~io26[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_1<=1001;io26[1:1]<=1;end
else if(m26_1<1250)begin m26_1<=m26_1+1;end
else if(m26_1==1250)begin m26_1<=0;io26[1:1]<=~io26[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_2<=407;io26[2:2]<=1;end
else if(m26_2<1250)begin m26_2<=m26_2+1;end
else if(m26_2==1250)begin m26_2<=0;io26[2:2]<=~io26[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_3<=493;io26[3:3]<=0;end
else if(m26_3<1250)begin m26_3<=m26_3+1;end
else if(m26_3==1250)begin m26_3<=0;io26[3:3]<=~io26[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_4<=164;io26[4:4]<=1;end
else if(m26_4<1250)begin m26_4<=m26_4+1;end
else if(m26_4==1250)begin m26_4<=0;io26[4:4]<=~io26[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_5<=648;io26[5:5]<=0;end
else if(m26_5<1250)begin m26_5<=m26_5+1;end
else if(m26_5==1250)begin m26_5<=0;io26[5:5]<=~io26[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_6<=719;io26[6:6]<=1;end
else if(m26_6<1250)begin m26_6<=m26_6+1;end
else if(m26_6==1250)begin m26_6<=0;io26[6:6]<=~io26[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_7<=534;io26[7:7]<=0;end
else if(m26_7<1250)begin m26_7<=m26_7+1;end
else if(m26_7==1250)begin m26_7<=0;io26[7:7]<=~io26[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_8<=1248;io26[8:8]<=0;end
else if(m26_8<1250)begin m26_8<=m26_8+1;end
else if(m26_8==1250)begin m26_8<=0;io26[8:8]<=~io26[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_9<=119;io26[9:9]<=1;end
else if(m26_9<1250)begin m26_9<=m26_9+1;end
else if(m26_9==1250)begin m26_9<=0;io26[9:9]<=~io26[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_10<=223;io26[10:10]<=0;end
else if(m26_10<1250)begin m26_10<=m26_10+1;end
else if(m26_10==1250)begin m26_10<=0;io26[10:10]<=~io26[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_11<=310;io26[11:11]<=0;end
else if(m26_11<1250)begin m26_11<=m26_11+1;end
else if(m26_11==1250)begin m26_11<=0;io26[11:11]<=~io26[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_12<=428;io26[12:12]<=0;end
else if(m26_12<1250)begin m26_12<=m26_12+1;end
else if(m26_12==1250)begin m26_12<=0;io26[12:12]<=~io26[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_13<=923;io26[13:13]<=1;end
else if(m26_13<1250)begin m26_13<=m26_13+1;end
else if(m26_13==1250)begin m26_13<=0;io26[13:13]<=~io26[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_14<=871;io26[14:14]<=0;end
else if(m26_14<1250)begin m26_14<=m26_14+1;end
else if(m26_14==1250)begin m26_14<=0;io26[14:14]<=~io26[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_15<=828;io26[15:15]<=0;end
else if(m26_15<1250)begin m26_15<=m26_15+1;end
else if(m26_15==1250)begin m26_15<=0;io26[15:15]<=~io26[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_16<=1154;io26[16:16]<=0;end
else if(m26_16<1250)begin m26_16<=m26_16+1;end
else if(m26_16==1250)begin m26_16<=0;io26[16:16]<=~io26[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_17<=910;io26[17:17]<=0;end
else if(m26_17<1250)begin m26_17<=m26_17+1;end
else if(m26_17==1250)begin m26_17<=0;io26[17:17]<=~io26[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_18<=336;io26[18:18]<=0;end
else if(m26_18<1250)begin m26_18<=m26_18+1;end
else if(m26_18==1250)begin m26_18<=0;io26[18:18]<=~io26[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_19<=237;io26[19:19]<=1;end
else if(m26_19<1250)begin m26_19<=m26_19+1;end
else if(m26_19==1250)begin m26_19<=0;io26[19:19]<=~io26[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_20<=1032;io26[20:20]<=1;end
else if(m26_20<1250)begin m26_20<=m26_20+1;end
else if(m26_20==1250)begin m26_20<=0;io26[20:20]<=~io26[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_21<=1112;io26[21:21]<=1;end
else if(m26_21<1250)begin m26_21<=m26_21+1;end
else if(m26_21==1250)begin m26_21<=0;io26[21:21]<=~io26[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_22<=1045;io26[22:22]<=1;end
else if(m26_22<1250)begin m26_22<=m26_22+1;end
else if(m26_22==1250)begin m26_22<=0;io26[22:22]<=~io26[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_23<=263;io26[23:23]<=1;end
else if(m26_23<1250)begin m26_23<=m26_23+1;end
else if(m26_23==1250)begin m26_23<=0;io26[23:23]<=~io26[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m26_24<=309;io26[24:24]<=0;end
else if(m26_24<1250)begin m26_24<=m26_24+1;end
else if(m26_24==1250)begin m26_24<=0;io26[24:24]<=~io26[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_0<=1084;io27[0:0]<=1;end
else if(m27_0<1250)begin m27_0<=m27_0+1;end
else if(m27_0==1250)begin m27_0<=0;io27[0:0]<=~io27[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_1<=1150;io27[1:1]<=1;end
else if(m27_1<1250)begin m27_1<=m27_1+1;end
else if(m27_1==1250)begin m27_1<=0;io27[1:1]<=~io27[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_2<=504;io27[2:2]<=1;end
else if(m27_2<1250)begin m27_2<=m27_2+1;end
else if(m27_2==1250)begin m27_2<=0;io27[2:2]<=~io27[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_3<=563;io27[3:3]<=0;end
else if(m27_3<1250)begin m27_3<=m27_3+1;end
else if(m27_3==1250)begin m27_3<=0;io27[3:3]<=~io27[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_4<=156;io27[4:4]<=1;end
else if(m27_4<1250)begin m27_4<=m27_4+1;end
else if(m27_4==1250)begin m27_4<=0;io27[4:4]<=~io27[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_5<=574;io27[5:5]<=0;end
else if(m27_5<1250)begin m27_5<=m27_5+1;end
else if(m27_5==1250)begin m27_5<=0;io27[5:5]<=~io27[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_6<=735;io27[6:6]<=1;end
else if(m27_6<1250)begin m27_6<=m27_6+1;end
else if(m27_6==1250)begin m27_6<=0;io27[6:6]<=~io27[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_7<=638;io27[7:7]<=0;end
else if(m27_7<1250)begin m27_7<=m27_7+1;end
else if(m27_7==1250)begin m27_7<=0;io27[7:7]<=~io27[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_8<=96;io27[8:8]<=1;end
else if(m27_8<1250)begin m27_8<=m27_8+1;end
else if(m27_8==1250)begin m27_8<=0;io27[8:8]<=~io27[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_9<=300;io27[9:9]<=1;end
else if(m27_9<1250)begin m27_9<=m27_9+1;end
else if(m27_9==1250)begin m27_9<=0;io27[9:9]<=~io27[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_10<=27;io27[10:10]<=0;end
else if(m27_10<1250)begin m27_10<=m27_10+1;end
else if(m27_10==1250)begin m27_10<=0;io27[10:10]<=~io27[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_11<=216;io27[11:11]<=0;end
else if(m27_11<1250)begin m27_11<=m27_11+1;end
else if(m27_11==1250)begin m27_11<=0;io27[11:11]<=~io27[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_12<=400;io27[12:12]<=0;end
else if(m27_12<1250)begin m27_12<=m27_12+1;end
else if(m27_12==1250)begin m27_12<=0;io27[12:12]<=~io27[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_13<=975;io27[13:13]<=1;end
else if(m27_13<1250)begin m27_13<=m27_13+1;end
else if(m27_13==1250)begin m27_13<=0;io27[13:13]<=~io27[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_14<=996;io27[14:14]<=0;end
else if(m27_14<1250)begin m27_14<=m27_14+1;end
else if(m27_14==1250)begin m27_14<=0;io27[14:14]<=~io27[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_15<=653;io27[15:15]<=0;end
else if(m27_15<1250)begin m27_15<=m27_15+1;end
else if(m27_15==1250)begin m27_15<=0;io27[15:15]<=~io27[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_16<=1005;io27[16:16]<=0;end
else if(m27_16<1250)begin m27_16<=m27_16+1;end
else if(m27_16==1250)begin m27_16<=0;io27[16:16]<=~io27[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_17<=855;io27[17:17]<=0;end
else if(m27_17<1250)begin m27_17<=m27_17+1;end
else if(m27_17==1250)begin m27_17<=0;io27[17:17]<=~io27[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_18<=292;io27[18:18]<=0;end
else if(m27_18<1250)begin m27_18<=m27_18+1;end
else if(m27_18==1250)begin m27_18<=0;io27[18:18]<=~io27[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_19<=275;io27[19:19]<=1;end
else if(m27_19<1250)begin m27_19<=m27_19+1;end
else if(m27_19==1250)begin m27_19<=0;io27[19:19]<=~io27[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_20<=827;io27[20:20]<=1;end
else if(m27_20<1250)begin m27_20<=m27_20+1;end
else if(m27_20==1250)begin m27_20<=0;io27[20:20]<=~io27[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_21<=944;io27[21:21]<=1;end
else if(m27_21<1250)begin m27_21<=m27_21+1;end
else if(m27_21==1250)begin m27_21<=0;io27[21:21]<=~io27[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_22<=894;io27[22:22]<=1;end
else if(m27_22<1250)begin m27_22<=m27_22+1;end
else if(m27_22==1250)begin m27_22<=0;io27[22:22]<=~io27[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_23<=216;io27[23:23]<=1;end
else if(m27_23<1250)begin m27_23<=m27_23+1;end
else if(m27_23==1250)begin m27_23<=0;io27[23:23]<=~io27[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m27_24<=283;io27[24:24]<=0;end
else if(m27_24<1250)begin m27_24<=m27_24+1;end
else if(m27_24==1250)begin m27_24<=0;io27[24:24]<=~io27[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_0<=1084;io28[0:0]<=1;end
else if(m28_0<1250)begin m28_0<=m28_0+1;end
else if(m28_0==1250)begin m28_0<=0;io28[0:0]<=~io28[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_1<=1150;io28[1:1]<=1;end
else if(m28_1<1250)begin m28_1<=m28_1+1;end
else if(m28_1==1250)begin m28_1<=0;io28[1:1]<=~io28[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_2<=504;io28[2:2]<=1;end
else if(m28_2<1250)begin m28_2<=m28_2+1;end
else if(m28_2==1250)begin m28_2<=0;io28[2:2]<=~io28[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_3<=563;io28[3:3]<=0;end
else if(m28_3<1250)begin m28_3<=m28_3+1;end
else if(m28_3==1250)begin m28_3<=0;io28[3:3]<=~io28[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_4<=156;io28[4:4]<=1;end
else if(m28_4<1250)begin m28_4<=m28_4+1;end
else if(m28_4==1250)begin m28_4<=0;io28[4:4]<=~io28[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_5<=574;io28[5:5]<=0;end
else if(m28_5<1250)begin m28_5<=m28_5+1;end
else if(m28_5==1250)begin m28_5<=0;io28[5:5]<=~io28[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_6<=735;io28[6:6]<=1;end
else if(m28_6<1250)begin m28_6<=m28_6+1;end
else if(m28_6==1250)begin m28_6<=0;io28[6:6]<=~io28[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_7<=638;io28[7:7]<=0;end
else if(m28_7<1250)begin m28_7<=m28_7+1;end
else if(m28_7==1250)begin m28_7<=0;io28[7:7]<=~io28[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_8<=96;io28[8:8]<=1;end
else if(m28_8<1250)begin m28_8<=m28_8+1;end
else if(m28_8==1250)begin m28_8<=0;io28[8:8]<=~io28[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_9<=300;io28[9:9]<=1;end
else if(m28_9<1250)begin m28_9<=m28_9+1;end
else if(m28_9==1250)begin m28_9<=0;io28[9:9]<=~io28[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_10<=27;io28[10:10]<=0;end
else if(m28_10<1250)begin m28_10<=m28_10+1;end
else if(m28_10==1250)begin m28_10<=0;io28[10:10]<=~io28[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_11<=216;io28[11:11]<=0;end
else if(m28_11<1250)begin m28_11<=m28_11+1;end
else if(m28_11==1250)begin m28_11<=0;io28[11:11]<=~io28[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_12<=400;io28[12:12]<=0;end
else if(m28_12<1250)begin m28_12<=m28_12+1;end
else if(m28_12==1250)begin m28_12<=0;io28[12:12]<=~io28[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_13<=975;io28[13:13]<=1;end
else if(m28_13<1250)begin m28_13<=m28_13+1;end
else if(m28_13==1250)begin m28_13<=0;io28[13:13]<=~io28[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_14<=996;io28[14:14]<=0;end
else if(m28_14<1250)begin m28_14<=m28_14+1;end
else if(m28_14==1250)begin m28_14<=0;io28[14:14]<=~io28[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_15<=653;io28[15:15]<=0;end
else if(m28_15<1250)begin m28_15<=m28_15+1;end
else if(m28_15==1250)begin m28_15<=0;io28[15:15]<=~io28[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_16<=1005;io28[16:16]<=0;end
else if(m28_16<1250)begin m28_16<=m28_16+1;end
else if(m28_16==1250)begin m28_16<=0;io28[16:16]<=~io28[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_17<=855;io28[17:17]<=0;end
else if(m28_17<1250)begin m28_17<=m28_17+1;end
else if(m28_17==1250)begin m28_17<=0;io28[17:17]<=~io28[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_18<=292;io28[18:18]<=0;end
else if(m28_18<1250)begin m28_18<=m28_18+1;end
else if(m28_18==1250)begin m28_18<=0;io28[18:18]<=~io28[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_19<=275;io28[19:19]<=1;end
else if(m28_19<1250)begin m28_19<=m28_19+1;end
else if(m28_19==1250)begin m28_19<=0;io28[19:19]<=~io28[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_20<=827;io28[20:20]<=1;end
else if(m28_20<1250)begin m28_20<=m28_20+1;end
else if(m28_20==1250)begin m28_20<=0;io28[20:20]<=~io28[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_21<=944;io28[21:21]<=1;end
else if(m28_21<1250)begin m28_21<=m28_21+1;end
else if(m28_21==1250)begin m28_21<=0;io28[21:21]<=~io28[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_22<=894;io28[22:22]<=1;end
else if(m28_22<1250)begin m28_22<=m28_22+1;end
else if(m28_22==1250)begin m28_22<=0;io28[22:22]<=~io28[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_23<=216;io28[23:23]<=1;end
else if(m28_23<1250)begin m28_23<=m28_23+1;end
else if(m28_23==1250)begin m28_23<=0;io28[23:23]<=~io28[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m28_24<=283;io28[24:24]<=0;end
else if(m28_24<1250)begin m28_24<=m28_24+1;end
else if(m28_24==1250)begin m28_24<=0;io28[24:24]<=~io28[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_0<=148;io29[0:0]<=0;end
else if(m29_0<1250)begin m29_0<=m29_0+1;end
else if(m29_0==1250)begin m29_0<=0;io29[0:0]<=~io29[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_1<=210;io29[1:1]<=0;end
else if(m29_1<1250)begin m29_1<=m29_1+1;end
else if(m29_1==1250)begin m29_1<=0;io29[1:1]<=~io29[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_2<=835;io29[2:2]<=1;end
else if(m29_2<1250)begin m29_2<=m29_2+1;end
else if(m29_2==1250)begin m29_2<=0;io29[2:2]<=~io29[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_3<=906;io29[3:3]<=0;end
else if(m29_3<1250)begin m29_3<=m29_3+1;end
else if(m29_3==1250)begin m29_3<=0;io29[3:3]<=~io29[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_4<=451;io29[4:4]<=1;end
else if(m29_4<1250)begin m29_4<=m29_4+1;end
else if(m29_4==1250)begin m29_4<=0;io29[4:4]<=~io29[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_5<=893;io29[5:5]<=0;end
else if(m29_5<1250)begin m29_5<=m29_5+1;end
else if(m29_5==1250)begin m29_5<=0;io29[5:5]<=~io29[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_6<=1010;io29[6:6]<=1;end
else if(m29_6<1250)begin m29_6<=m29_6+1;end
else if(m29_6==1250)begin m29_6<=0;io29[6:6]<=~io29[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_7<=913;io29[7:7]<=0;end
else if(m29_7<1250)begin m29_7<=m29_7+1;end
else if(m29_7==1250)begin m29_7<=0;io29[7:7]<=~io29[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_8<=362;io29[8:8]<=1;end
else if(m29_8<1250)begin m29_8<=m29_8+1;end
else if(m29_8==1250)begin m29_8<=0;io29[8:8]<=~io29[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_9<=555;io29[9:9]<=1;end
else if(m29_9<1250)begin m29_9<=m29_9+1;end
else if(m29_9==1250)begin m29_9<=0;io29[9:9]<=~io29[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_10<=202;io29[10:10]<=0;end
else if(m29_10<1250)begin m29_10<=m29_10+1;end
else if(m29_10==1250)begin m29_10<=0;io29[10:10]<=~io29[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_11<=390;io29[11:11]<=0;end
else if(m29_11<1250)begin m29_11<=m29_11+1;end
else if(m29_11==1250)begin m29_11<=0;io29[11:11]<=~io29[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_12<=570;io29[12:12]<=0;end
else if(m29_12<1250)begin m29_12<=m29_12+1;end
else if(m29_12==1250)begin m29_12<=0;io29[12:12]<=~io29[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_13<=1162;io29[13:13]<=1;end
else if(m29_13<1250)begin m29_13<=m29_13+1;end
else if(m29_13==1250)begin m29_13<=0;io29[13:13]<=~io29[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_14<=1185;io29[14:14]<=0;end
else if(m29_14<1250)begin m29_14<=m29_14+1;end
else if(m29_14==1250)begin m29_14<=0;io29[14:14]<=~io29[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_15<=752;io29[15:15]<=0;end
else if(m29_15<1250)begin m29_15<=m29_15+1;end
else if(m29_15==1250)begin m29_15<=0;io29[15:15]<=~io29[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_16<=1126;io29[16:16]<=0;end
else if(m29_16<1250)begin m29_16<=m29_16+1;end
else if(m29_16==1250)begin m29_16<=0;io29[16:16]<=~io29[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_17<=986;io29[17:17]<=0;end
else if(m29_17<1250)begin m29_17<=m29_17+1;end
else if(m29_17==1250)begin m29_17<=0;io29[17:17]<=~io29[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_18<=393;io29[18:18]<=0;end
else if(m29_18<1250)begin m29_18<=m29_18+1;end
else if(m29_18==1250)begin m29_18<=0;io29[18:18]<=~io29[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_19<=406;io29[19:19]<=1;end
else if(m29_19<1250)begin m29_19<=m29_19+1;end
else if(m29_19==1250)begin m29_19<=0;io29[19:19]<=~io29[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_20<=803;io29[20:20]<=1;end
else if(m29_20<1250)begin m29_20<=m29_20+1;end
else if(m29_20==1250)begin m29_20<=0;io29[20:20]<=~io29[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_21<=1022;io29[21:21]<=1;end
else if(m29_21<1250)begin m29_21<=m29_21+1;end
else if(m29_21==1250)begin m29_21<=0;io29[21:21]<=~io29[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_22<=954;io29[22:22]<=1;end
else if(m29_22<1250)begin m29_22<=m29_22+1;end
else if(m29_22==1250)begin m29_22<=0;io29[22:22]<=~io29[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_23<=223;io29[23:23]<=1;end
else if(m29_23<1250)begin m29_23<=m29_23+1;end
else if(m29_23==1250)begin m29_23<=0;io29[23:23]<=~io29[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m29_24<=360;io29[24:24]<=0;end
else if(m29_24<1250)begin m29_24<=m29_24+1;end
else if(m29_24==1250)begin m29_24<=0;io29[24:24]<=~io29[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_0<=269;io30[0:0]<=0;end
else if(m30_0<1250)begin m30_0<=m30_0+1;end
else if(m30_0==1250)begin m30_0<=0;io30[0:0]<=~io30[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_1<=361;io30[1:1]<=0;end
else if(m30_1<1250)begin m30_1<=m30_1+1;end
else if(m30_1==1250)begin m30_1<=0;io30[1:1]<=~io30[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_2<=981;io30[2:2]<=1;end
else if(m30_2<1250)begin m30_2<=m30_2+1;end
else if(m30_2==1250)begin m30_2<=0;io30[2:2]<=~io30[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_3<=1043;io30[3:3]<=0;end
else if(m30_3<1250)begin m30_3<=m30_3+1;end
else if(m30_3==1250)begin m30_3<=0;io30[3:3]<=~io30[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_4<=623;io30[4:4]<=1;end
else if(m30_4<1250)begin m30_4<=m30_4+1;end
else if(m30_4==1250)begin m30_4<=0;io30[4:4]<=~io30[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_5<=1023;io30[5:5]<=0;end
else if(m30_5<1250)begin m30_5<=m30_5+1;end
else if(m30_5==1250)begin m30_5<=0;io30[5:5]<=~io30[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_6<=1085;io30[6:6]<=1;end
else if(m30_6<1250)begin m30_6<=m30_6+1;end
else if(m30_6==1250)begin m30_6<=0;io30[6:6]<=~io30[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_7<=986;io30[7:7]<=0;end
else if(m30_7<1250)begin m30_7<=m30_7+1;end
else if(m30_7==1250)begin m30_7<=0;io30[7:7]<=~io30[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_8<=456;io30[8:8]<=1;end
else if(m30_8<1250)begin m30_8<=m30_8+1;end
else if(m30_8==1250)begin m30_8<=0;io30[8:8]<=~io30[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_9<=615;io30[9:9]<=1;end
else if(m30_9<1250)begin m30_9<=m30_9+1;end
else if(m30_9==1250)begin m30_9<=0;io30[9:9]<=~io30[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_10<=202;io30[10:10]<=0;end
else if(m30_10<1250)begin m30_10<=m30_10+1;end
else if(m30_10==1250)begin m30_10<=0;io30[10:10]<=~io30[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_11<=390;io30[11:11]<=0;end
else if(m30_11<1250)begin m30_11<=m30_11+1;end
else if(m30_11==1250)begin m30_11<=0;io30[11:11]<=~io30[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_12<=570;io30[12:12]<=0;end
else if(m30_12<1250)begin m30_12<=m30_12+1;end
else if(m30_12==1250)begin m30_12<=0;io30[12:12]<=~io30[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_13<=1162;io30[13:13]<=1;end
else if(m30_13<1250)begin m30_13<=m30_13+1;end
else if(m30_13==1250)begin m30_13<=0;io30[13:13]<=~io30[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_14<=1185;io30[14:14]<=0;end
else if(m30_14<1250)begin m30_14<=m30_14+1;end
else if(m30_14==1250)begin m30_14<=0;io30[14:14]<=~io30[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_15<=622;io30[15:15]<=0;end
else if(m30_15<1250)begin m30_15<=m30_15+1;end
else if(m30_15==1250)begin m30_15<=0;io30[15:15]<=~io30[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_16<=1052;io30[16:16]<=0;end
else if(m30_16<1250)begin m30_16<=m30_16+1;end
else if(m30_16==1250)begin m30_16<=0;io30[16:16]<=~io30[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_17<=913;io30[17:17]<=0;end
else if(m30_17<1250)begin m30_17<=m30_17+1;end
else if(m30_17==1250)begin m30_17<=0;io30[17:17]<=~io30[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_18<=299;io30[18:18]<=0;end
else if(m30_18<1250)begin m30_18<=m30_18+1;end
else if(m30_18==1250)begin m30_18<=0;io30[18:18]<=~io30[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_19<=346;io30[19:19]<=1;end
else if(m30_19<1250)begin m30_19<=m30_19+1;end
else if(m30_19==1250)begin m30_19<=0;io30[19:19]<=~io30[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_20<=632;io30[20:20]<=1;end
else if(m30_20<1250)begin m30_20<=m30_20+1;end
else if(m30_20==1250)begin m30_20<=0;io30[20:20]<=~io30[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_21<=885;io30[21:21]<=1;end
else if(m30_21<1250)begin m30_21<=m30_21+1;end
else if(m30_21==1250)begin m30_21<=0;io30[21:21]<=~io30[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_22<=808;io30[22:22]<=1;end
else if(m30_22<1250)begin m30_22<=m30_22+1;end
else if(m30_22==1250)begin m30_22<=0;io30[22:22]<=~io30[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_23<=71;io30[23:23]<=1;end
else if(m30_23<1250)begin m30_23<=m30_23+1;end
else if(m30_23==1250)begin m30_23<=0;io30[23:23]<=~io30[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m30_24<=238;io30[24:24]<=0;end
else if(m30_24<1250)begin m30_24<=m30_24+1;end
else if(m30_24==1250)begin m30_24<=0;io30[24:24]<=~io30[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_0<=269;io31[0:0]<=0;end
else if(m31_0<1250)begin m31_0<=m31_0+1;end
else if(m31_0==1250)begin m31_0<=0;io31[0:0]<=~io31[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_1<=361;io31[1:1]<=0;end
else if(m31_1<1250)begin m31_1<=m31_1+1;end
else if(m31_1==1250)begin m31_1<=0;io31[1:1]<=~io31[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_2<=981;io31[2:2]<=1;end
else if(m31_2<1250)begin m31_2<=m31_2+1;end
else if(m31_2==1250)begin m31_2<=0;io31[2:2]<=~io31[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_3<=1043;io31[3:3]<=0;end
else if(m31_3<1250)begin m31_3<=m31_3+1;end
else if(m31_3==1250)begin m31_3<=0;io31[3:3]<=~io31[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_4<=623;io31[4:4]<=1;end
else if(m31_4<1250)begin m31_4<=m31_4+1;end
else if(m31_4==1250)begin m31_4<=0;io31[4:4]<=~io31[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_5<=1023;io31[5:5]<=0;end
else if(m31_5<1250)begin m31_5<=m31_5+1;end
else if(m31_5==1250)begin m31_5<=0;io31[5:5]<=~io31[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_6<=1085;io31[6:6]<=1;end
else if(m31_6<1250)begin m31_6<=m31_6+1;end
else if(m31_6==1250)begin m31_6<=0;io31[6:6]<=~io31[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_7<=986;io31[7:7]<=0;end
else if(m31_7<1250)begin m31_7<=m31_7+1;end
else if(m31_7==1250)begin m31_7<=0;io31[7:7]<=~io31[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_8<=456;io31[8:8]<=1;end
else if(m31_8<1250)begin m31_8<=m31_8+1;end
else if(m31_8==1250)begin m31_8<=0;io31[8:8]<=~io31[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_9<=615;io31[9:9]<=1;end
else if(m31_9<1250)begin m31_9<=m31_9+1;end
else if(m31_9==1250)begin m31_9<=0;io31[9:9]<=~io31[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_10<=202;io31[10:10]<=0;end
else if(m31_10<1250)begin m31_10<=m31_10+1;end
else if(m31_10==1250)begin m31_10<=0;io31[10:10]<=~io31[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_11<=390;io31[11:11]<=0;end
else if(m31_11<1250)begin m31_11<=m31_11+1;end
else if(m31_11==1250)begin m31_11<=0;io31[11:11]<=~io31[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_12<=570;io31[12:12]<=0;end
else if(m31_12<1250)begin m31_12<=m31_12+1;end
else if(m31_12==1250)begin m31_12<=0;io31[12:12]<=~io31[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_13<=1162;io31[13:13]<=1;end
else if(m31_13<1250)begin m31_13<=m31_13+1;end
else if(m31_13==1250)begin m31_13<=0;io31[13:13]<=~io31[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_14<=1185;io31[14:14]<=0;end
else if(m31_14<1250)begin m31_14<=m31_14+1;end
else if(m31_14==1250)begin m31_14<=0;io31[14:14]<=~io31[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_15<=622;io31[15:15]<=0;end
else if(m31_15<1250)begin m31_15<=m31_15+1;end
else if(m31_15==1250)begin m31_15<=0;io31[15:15]<=~io31[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_16<=1052;io31[16:16]<=0;end
else if(m31_16<1250)begin m31_16<=m31_16+1;end
else if(m31_16==1250)begin m31_16<=0;io31[16:16]<=~io31[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_17<=913;io31[17:17]<=0;end
else if(m31_17<1250)begin m31_17<=m31_17+1;end
else if(m31_17==1250)begin m31_17<=0;io31[17:17]<=~io31[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_18<=299;io31[18:18]<=0;end
else if(m31_18<1250)begin m31_18<=m31_18+1;end
else if(m31_18==1250)begin m31_18<=0;io31[18:18]<=~io31[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_19<=346;io31[19:19]<=1;end
else if(m31_19<1250)begin m31_19<=m31_19+1;end
else if(m31_19==1250)begin m31_19<=0;io31[19:19]<=~io31[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_20<=632;io31[20:20]<=1;end
else if(m31_20<1250)begin m31_20<=m31_20+1;end
else if(m31_20==1250)begin m31_20<=0;io31[20:20]<=~io31[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_21<=885;io31[21:21]<=1;end
else if(m31_21<1250)begin m31_21<=m31_21+1;end
else if(m31_21==1250)begin m31_21<=0;io31[21:21]<=~io31[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_22<=808;io31[22:22]<=1;end
else if(m31_22<1250)begin m31_22<=m31_22+1;end
else if(m31_22==1250)begin m31_22<=0;io31[22:22]<=~io31[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_23<=71;io31[23:23]<=1;end
else if(m31_23<1250)begin m31_23<=m31_23+1;end
else if(m31_23==1250)begin m31_23<=0;io31[23:23]<=~io31[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m31_24<=238;io31[24:24]<=0;end
else if(m31_24<1250)begin m31_24<=m31_24+1;end
else if(m31_24==1250)begin m31_24<=0;io31[24:24]<=~io31[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_0<=348;io32[0:0]<=0;end
else if(m32_0<1250)begin m32_0<=m32_0+1;end
else if(m32_0==1250)begin m32_0<=0;io32[0:0]<=~io32[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_1<=522;io32[1:1]<=0;end
else if(m32_1<1250)begin m32_1<=m32_1+1;end
else if(m32_1==1250)begin m32_1<=0;io32[1:1]<=~io32[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_2<=1197;io32[2:2]<=1;end
else if(m32_2<1250)begin m32_2<=m32_2+1;end
else if(m32_2==1250)begin m32_2<=0;io32[2:2]<=~io32[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_3<=23;io32[3:3]<=1;end
else if(m32_3<1250)begin m32_3<=m32_3+1;end
else if(m32_3==1250)begin m32_3<=0;io32[3:3]<=~io32[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_4<=955;io32[4:4]<=1;end
else if(m32_4<1250)begin m32_4<=m32_4+1;end
else if(m32_4==1250)begin m32_4<=0;io32[4:4]<=~io32[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_5<=52;io32[5:5]<=1;end
else if(m32_5<1250)begin m32_5<=m32_5+1;end
else if(m32_5==1250)begin m32_5<=0;io32[5:5]<=~io32[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_6<=30;io32[6:6]<=0;end
else if(m32_6<1250)begin m32_6<=m32_6+1;end
else if(m32_6==1250)begin m32_6<=0;io32[6:6]<=~io32[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_7<=1098;io32[7:7]<=0;end
else if(m32_7<1250)begin m32_7<=m32_7+1;end
else if(m32_7==1250)begin m32_7<=0;io32[7:7]<=~io32[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_8<=570;io32[8:8]<=1;end
else if(m32_8<1250)begin m32_8<=m32_8+1;end
else if(m32_8==1250)begin m32_8<=0;io32[8:8]<=~io32[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_9<=635;io32[9:9]<=1;end
else if(m32_9<1250)begin m32_9<=m32_9+1;end
else if(m32_9==1250)begin m32_9<=0;io32[9:9]<=~io32[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_10<=416;io32[10:10]<=0;end
else if(m32_10<1250)begin m32_10<=m32_10+1;end
else if(m32_10==1250)begin m32_10<=0;io32[10:10]<=~io32[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_11<=529;io32[11:11]<=0;end
else if(m32_11<1250)begin m32_11<=m32_11+1;end
else if(m32_11==1250)begin m32_11<=0;io32[11:11]<=~io32[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_12<=636;io32[12:12]<=0;end
else if(m32_12<1250)begin m32_12<=m32_12+1;end
else if(m32_12==1250)begin m32_12<=0;io32[12:12]<=~io32[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_13<=1159;io32[13:13]<=1;end
else if(m32_13<1250)begin m32_13<=m32_13+1;end
else if(m32_13==1250)begin m32_13<=0;io32[13:13]<=~io32[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_14<=1114;io32[14:14]<=0;end
else if(m32_14<1250)begin m32_14<=m32_14+1;end
else if(m32_14==1250)begin m32_14<=0;io32[14:14]<=~io32[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_15<=717;io32[15:15]<=0;end
else if(m32_15<1250)begin m32_15<=m32_15+1;end
else if(m32_15==1250)begin m32_15<=0;io32[15:15]<=~io32[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_16<=1093;io32[16:16]<=0;end
else if(m32_16<1250)begin m32_16<=m32_16+1;end
else if(m32_16==1250)begin m32_16<=0;io32[16:16]<=~io32[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_17<=865;io32[17:17]<=0;end
else if(m32_17<1250)begin m32_17<=m32_17+1;end
else if(m32_17==1250)begin m32_17<=0;io32[17:17]<=~io32[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_18<=234;io32[18:18]<=0;end
else if(m32_18<1250)begin m32_18<=m32_18+1;end
else if(m32_18==1250)begin m32_18<=0;io32[18:18]<=~io32[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_19<=235;io32[19:19]<=1;end
else if(m32_19<1250)begin m32_19<=m32_19+1;end
else if(m32_19==1250)begin m32_19<=0;io32[19:19]<=~io32[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_20<=661;io32[20:20]<=1;end
else if(m32_20<1250)begin m32_20<=m32_20+1;end
else if(m32_20==1250)begin m32_20<=0;io32[20:20]<=~io32[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_21<=861;io32[21:21]<=1;end
else if(m32_21<1250)begin m32_21<=m32_21+1;end
else if(m32_21==1250)begin m32_21<=0;io32[21:21]<=~io32[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_22<=745;io32[22:22]<=1;end
else if(m32_22<1250)begin m32_22<=m32_22+1;end
else if(m32_22==1250)begin m32_22<=0;io32[22:22]<=~io32[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_23<=1225;io32[23:23]<=0;end
else if(m32_23<1250)begin m32_23<=m32_23+1;end
else if(m32_23==1250)begin m32_23<=0;io32[23:23]<=~io32[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m32_24<=91;io32[24:24]<=0;end
else if(m32_24<1250)begin m32_24<=m32_24+1;end
else if(m32_24==1250)begin m32_24<=0;io32[24:24]<=~io32[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_0<=348;io33[0:0]<=0;end
else if(m33_0<1250)begin m33_0<=m33_0+1;end
else if(m33_0==1250)begin m33_0<=0;io33[0:0]<=~io33[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_1<=522;io33[1:1]<=0;end
else if(m33_1<1250)begin m33_1<=m33_1+1;end
else if(m33_1==1250)begin m33_1<=0;io33[1:1]<=~io33[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_2<=1197;io33[2:2]<=1;end
else if(m33_2<1250)begin m33_2<=m33_2+1;end
else if(m33_2==1250)begin m33_2<=0;io33[2:2]<=~io33[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_3<=23;io33[3:3]<=1;end
else if(m33_3<1250)begin m33_3<=m33_3+1;end
else if(m33_3==1250)begin m33_3<=0;io33[3:3]<=~io33[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_4<=955;io33[4:4]<=1;end
else if(m33_4<1250)begin m33_4<=m33_4+1;end
else if(m33_4==1250)begin m33_4<=0;io33[4:4]<=~io33[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_5<=52;io33[5:5]<=1;end
else if(m33_5<1250)begin m33_5<=m33_5+1;end
else if(m33_5==1250)begin m33_5<=0;io33[5:5]<=~io33[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_6<=30;io33[6:6]<=0;end
else if(m33_6<1250)begin m33_6<=m33_6+1;end
else if(m33_6==1250)begin m33_6<=0;io33[6:6]<=~io33[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_7<=1098;io33[7:7]<=0;end
else if(m33_7<1250)begin m33_7<=m33_7+1;end
else if(m33_7==1250)begin m33_7<=0;io33[7:7]<=~io33[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_8<=570;io33[8:8]<=1;end
else if(m33_8<1250)begin m33_8<=m33_8+1;end
else if(m33_8==1250)begin m33_8<=0;io33[8:8]<=~io33[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_9<=635;io33[9:9]<=1;end
else if(m33_9<1250)begin m33_9<=m33_9+1;end
else if(m33_9==1250)begin m33_9<=0;io33[9:9]<=~io33[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_10<=416;io33[10:10]<=0;end
else if(m33_10<1250)begin m33_10<=m33_10+1;end
else if(m33_10==1250)begin m33_10<=0;io33[10:10]<=~io33[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_11<=529;io33[11:11]<=0;end
else if(m33_11<1250)begin m33_11<=m33_11+1;end
else if(m33_11==1250)begin m33_11<=0;io33[11:11]<=~io33[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_12<=636;io33[12:12]<=0;end
else if(m33_12<1250)begin m33_12<=m33_12+1;end
else if(m33_12==1250)begin m33_12<=0;io33[12:12]<=~io33[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_13<=1159;io33[13:13]<=1;end
else if(m33_13<1250)begin m33_13<=m33_13+1;end
else if(m33_13==1250)begin m33_13<=0;io33[13:13]<=~io33[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_14<=1114;io33[14:14]<=0;end
else if(m33_14<1250)begin m33_14<=m33_14+1;end
else if(m33_14==1250)begin m33_14<=0;io33[14:14]<=~io33[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_15<=717;io33[15:15]<=0;end
else if(m33_15<1250)begin m33_15<=m33_15+1;end
else if(m33_15==1250)begin m33_15<=0;io33[15:15]<=~io33[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_16<=1093;io33[16:16]<=0;end
else if(m33_16<1250)begin m33_16<=m33_16+1;end
else if(m33_16==1250)begin m33_16<=0;io33[16:16]<=~io33[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_17<=865;io33[17:17]<=0;end
else if(m33_17<1250)begin m33_17<=m33_17+1;end
else if(m33_17==1250)begin m33_17<=0;io33[17:17]<=~io33[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_18<=234;io33[18:18]<=0;end
else if(m33_18<1250)begin m33_18<=m33_18+1;end
else if(m33_18==1250)begin m33_18<=0;io33[18:18]<=~io33[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_19<=235;io33[19:19]<=1;end
else if(m33_19<1250)begin m33_19<=m33_19+1;end
else if(m33_19==1250)begin m33_19<=0;io33[19:19]<=~io33[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_20<=661;io33[20:20]<=1;end
else if(m33_20<1250)begin m33_20<=m33_20+1;end
else if(m33_20==1250)begin m33_20<=0;io33[20:20]<=~io33[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_21<=861;io33[21:21]<=1;end
else if(m33_21<1250)begin m33_21<=m33_21+1;end
else if(m33_21==1250)begin m33_21<=0;io33[21:21]<=~io33[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_22<=745;io33[22:22]<=1;end
else if(m33_22<1250)begin m33_22<=m33_22+1;end
else if(m33_22==1250)begin m33_22<=0;io33[22:22]<=~io33[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_23<=1225;io33[23:23]<=0;end
else if(m33_23<1250)begin m33_23<=m33_23+1;end
else if(m33_23==1250)begin m33_23<=0;io33[23:23]<=~io33[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m33_24<=91;io33[24:24]<=0;end
else if(m33_24<1250)begin m33_24<=m33_24+1;end
else if(m33_24==1250)begin m33_24<=0;io33[24:24]<=~io33[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_0<=219;io34[0:0]<=0;end
else if(m34_0<1250)begin m34_0<=m34_0+1;end
else if(m34_0==1250)begin m34_0<=0;io34[0:0]<=~io34[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_1<=402;io34[1:1]<=0;end
else if(m34_1<1250)begin m34_1<=m34_1+1;end
else if(m34_1==1250)begin m34_1<=0;io34[1:1]<=~io34[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_2<=1073;io34[2:2]<=1;end
else if(m34_2<1250)begin m34_2<=m34_2+1;end
else if(m34_2==1250)begin m34_2<=0;io34[2:2]<=~io34[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_3<=1132;io34[3:3]<=0;end
else if(m34_3<1250)begin m34_3<=m34_3+1;end
else if(m34_3==1250)begin m34_3<=0;io34[3:3]<=~io34[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_4<=852;io34[4:4]<=1;end
else if(m34_4<1250)begin m34_4<=m34_4+1;end
else if(m34_4==1250)begin m34_4<=0;io34[4:4]<=~io34[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_5<=1099;io34[5:5]<=0;end
else if(m34_5<1250)begin m34_5<=m34_5+1;end
else if(m34_5==1250)begin m34_5<=0;io34[5:5]<=~io34[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_6<=1112;io34[6:6]<=1;end
else if(m34_6<1250)begin m34_6<=m34_6+1;end
else if(m34_6==1250)begin m34_6<=0;io34[6:6]<=~io34[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_7<=910;io34[7:7]<=0;end
else if(m34_7<1250)begin m34_7<=m34_7+1;end
else if(m34_7==1250)begin m34_7<=0;io34[7:7]<=~io34[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_8<=398;io34[8:8]<=1;end
else if(m34_8<1250)begin m34_8<=m34_8+1;end
else if(m34_8==1250)begin m34_8<=0;io34[8:8]<=~io34[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_9<=445;io34[9:9]<=1;end
else if(m34_9<1250)begin m34_9<=m34_9+1;end
else if(m34_9==1250)begin m34_9<=0;io34[9:9]<=~io34[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_10<=223;io34[10:10]<=0;end
else if(m34_10<1250)begin m34_10<=m34_10+1;end
else if(m34_10==1250)begin m34_10<=0;io34[10:10]<=~io34[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_11<=310;io34[11:11]<=0;end
else if(m34_11<1250)begin m34_11<=m34_11+1;end
else if(m34_11==1250)begin m34_11<=0;io34[11:11]<=~io34[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_12<=428;io34[12:12]<=0;end
else if(m34_12<1250)begin m34_12<=m34_12+1;end
else if(m34_12==1250)begin m34_12<=0;io34[12:12]<=~io34[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_13<=923;io34[13:13]<=1;end
else if(m34_13<1250)begin m34_13<=m34_13+1;end
else if(m34_13==1250)begin m34_13<=0;io34[13:13]<=~io34[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_14<=871;io34[14:14]<=0;end
else if(m34_14<1250)begin m34_14<=m34_14+1;end
else if(m34_14==1250)begin m34_14<=0;io34[14:14]<=~io34[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_15<=377;io34[15:15]<=0;end
else if(m34_15<1250)begin m34_15<=m34_15+1;end
else if(m34_15==1250)begin m34_15<=0;io34[15:15]<=~io34[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_16<=761;io34[16:16]<=0;end
else if(m34_16<1250)begin m34_16<=m34_16+1;end
else if(m34_16==1250)begin m34_16<=0;io34[16:16]<=~io34[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_17<=534;io34[17:17]<=0;end
else if(m34_17<1250)begin m34_17<=m34_17+1;end
else if(m34_17==1250)begin m34_17<=0;io34[17:17]<=~io34[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_18<=1186;io34[18:18]<=1;end
else if(m34_18<1250)begin m34_18<=m34_18+1;end
else if(m34_18==1250)begin m34_18<=0;io34[18:18]<=~io34[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_19<=1161;io34[19:19]<=0;end
else if(m34_19<1250)begin m34_19<=m34_19+1;end
else if(m34_19==1250)begin m34_19<=0;io34[19:19]<=~io34[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_20<=345;io34[20:20]<=1;end
else if(m34_20<1250)begin m34_20<=m34_20+1;end
else if(m34_20==1250)begin m34_20<=0;io34[20:20]<=~io34[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_21<=473;io34[21:21]<=1;end
else if(m34_21<1250)begin m34_21<=m34_21+1;end
else if(m34_21==1250)begin m34_21<=0;io34[21:21]<=~io34[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_22<=379;io34[22:22]<=1;end
else if(m34_22<1250)begin m34_22<=m34_22+1;end
else if(m34_22==1250)begin m34_22<=0;io34[22:22]<=~io34[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_23<=862;io34[23:23]<=0;end
else if(m34_23<1250)begin m34_23<=m34_23+1;end
else if(m34_23==1250)begin m34_23<=0;io34[23:23]<=~io34[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m34_24<=986;io34[24:24]<=1;end
else if(m34_24<1250)begin m34_24<=m34_24+1;end
else if(m34_24==1250)begin m34_24<=0;io34[24:24]<=~io34[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_0<=1233;io35[0:0]<=1;end
else if(m35_0<1250)begin m35_0<=m35_0+1;end
else if(m35_0==1250)begin m35_0<=0;io35[0:0]<=~io35[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_1<=178;io35[1:1]<=0;end
else if(m35_1<1250)begin m35_1<=m35_1+1;end
else if(m35_1==1250)begin m35_1<=0;io35[1:1]<=~io35[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_2<=970;io35[2:2]<=1;end
else if(m35_2<1250)begin m35_2<=m35_2+1;end
else if(m35_2==1250)begin m35_2<=0;io35[2:2]<=~io35[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_3<=1034;io35[3:3]<=0;end
else if(m35_3<1250)begin m35_3<=m35_3+1;end
else if(m35_3==1250)begin m35_3<=0;io35[3:3]<=~io35[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_4<=805;io35[4:4]<=1;end
else if(m35_4<1250)begin m35_4<=m35_4+1;end
else if(m35_4==1250)begin m35_4<=0;io35[4:4]<=~io35[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_5<=1045;io35[5:5]<=0;end
else if(m35_5<1250)begin m35_5<=m35_5+1;end
else if(m35_5==1250)begin m35_5<=0;io35[5:5]<=~io35[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_6<=1041;io35[6:6]<=1;end
else if(m35_6<1250)begin m35_6<=m35_6+1;end
else if(m35_6==1250)begin m35_6<=0;io35[6:6]<=~io35[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_7<=758;io35[7:7]<=0;end
else if(m35_7<1250)begin m35_7<=m35_7+1;end
else if(m35_7==1250)begin m35_7<=0;io35[7:7]<=~io35[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_8<=219;io35[8:8]<=1;end
else if(m35_8<1250)begin m35_8<=m35_8+1;end
else if(m35_8==1250)begin m35_8<=0;io35[8:8]<=~io35[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_9<=170;io35[9:9]<=1;end
else if(m35_9<1250)begin m35_9<=m35_9+1;end
else if(m35_9==1250)begin m35_9<=0;io35[9:9]<=~io35[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_10<=208;io35[10:10]<=0;end
else if(m35_10<1250)begin m35_10<=m35_10+1;end
else if(m35_10==1250)begin m35_10<=0;io35[10:10]<=~io35[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_11<=245;io35[11:11]<=0;end
else if(m35_11<1250)begin m35_11<=m35_11+1;end
else if(m35_11==1250)begin m35_11<=0;io35[11:11]<=~io35[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_12<=272;io35[12:12]<=0;end
else if(m35_12<1250)begin m35_12<=m35_12+1;end
else if(m35_12==1250)begin m35_12<=0;io35[12:12]<=~io35[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_13<=705;io35[13:13]<=1;end
else if(m35_13<1250)begin m35_13<=m35_13+1;end
else if(m35_13==1250)begin m35_13<=0;io35[13:13]<=~io35[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_14<=585;io35[14:14]<=0;end
else if(m35_14<1250)begin m35_14<=m35_14+1;end
else if(m35_14==1250)begin m35_14<=0;io35[14:14]<=~io35[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_15<=371;io35[15:15]<=0;end
else if(m35_15<1250)begin m35_15<=m35_15+1;end
else if(m35_15==1250)begin m35_15<=0;io35[15:15]<=~io35[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_16<=712;io35[16:16]<=0;end
else if(m35_16<1250)begin m35_16<=m35_16+1;end
else if(m35_16==1250)begin m35_16<=0;io35[16:16]<=~io35[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_17<=363;io35[17:17]<=0;end
else if(m35_17<1250)begin m35_17<=m35_17+1;end
else if(m35_17==1250)begin m35_17<=0;io35[17:17]<=~io35[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_18<=982;io35[18:18]<=1;end
else if(m35_18<1250)begin m35_18<=m35_18+1;end
else if(m35_18==1250)begin m35_18<=0;io35[18:18]<=~io35[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_19<=877;io35[19:19]<=0;end
else if(m35_19<1250)begin m35_19<=m35_19+1;end
else if(m35_19==1250)begin m35_19<=0;io35[19:19]<=~io35[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_20<=284;io35[20:20]<=1;end
else if(m35_20<1250)begin m35_20<=m35_20+1;end
else if(m35_20==1250)begin m35_20<=0;io35[20:20]<=~io35[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_21<=375;io35[21:21]<=1;end
else if(m35_21<1250)begin m35_21<=m35_21+1;end
else if(m35_21==1250)begin m35_21<=0;io35[21:21]<=~io35[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_22<=259;io35[22:22]<=1;end
else if(m35_22<1250)begin m35_22<=m35_22+1;end
else if(m35_22==1250)begin m35_22<=0;io35[22:22]<=~io35[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_23<=685;io35[23:23]<=0;end
else if(m35_23<1250)begin m35_23<=m35_23+1;end
else if(m35_23==1250)begin m35_23<=0;io35[23:23]<=~io35[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m35_24<=757;io35[24:24]<=1;end
else if(m35_24<1250)begin m35_24<=m35_24+1;end
else if(m35_24==1250)begin m35_24<=0;io35[24:24]<=~io35[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_0<=1052;io36[0:0]<=1;end
else if(m36_0<1250)begin m36_0<=m36_0+1;end
else if(m36_0==1250)begin m36_0<=0;io36[0:0]<=~io36[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_1<=1239;io36[1:1]<=1;end
else if(m36_1<1250)begin m36_1<=m36_1+1;end
else if(m36_1==1250)begin m36_1<=0;io36[1:1]<=~io36[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_2<=927;io36[2:2]<=1;end
else if(m36_2<1250)begin m36_2<=m36_2+1;end
else if(m36_2==1250)begin m36_2<=0;io36[2:2]<=~io36[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_3<=1006;io36[3:3]<=0;end
else if(m36_3<1250)begin m36_3<=m36_3+1;end
else if(m36_3==1250)begin m36_3<=0;io36[3:3]<=~io36[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_4<=849;io36[4:4]<=1;end
else if(m36_4<1250)begin m36_4<=m36_4+1;end
else if(m36_4==1250)begin m36_4<=0;io36[4:4]<=~io36[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_5<=959;io36[5:5]<=0;end
else if(m36_5<1250)begin m36_5<=m36_5+1;end
else if(m36_5==1250)begin m36_5<=0;io36[5:5]<=~io36[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_6<=985;io36[6:6]<=1;end
else if(m36_6<1250)begin m36_6<=m36_6+1;end
else if(m36_6==1250)begin m36_6<=0;io36[6:6]<=~io36[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_7<=624;io36[7:7]<=0;end
else if(m36_7<1250)begin m36_7<=m36_7+1;end
else if(m36_7==1250)begin m36_7<=0;io36[7:7]<=~io36[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_8<=19;io36[8:8]<=1;end
else if(m36_8<1250)begin m36_8<=m36_8+1;end
else if(m36_8==1250)begin m36_8<=0;io36[8:8]<=~io36[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_9<=1138;io36[9:9]<=0;end
else if(m36_9<1250)begin m36_9<=m36_9+1;end
else if(m36_9==1250)begin m36_9<=0;io36[9:9]<=~io36[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_10<=187;io36[10:10]<=0;end
else if(m36_10<1250)begin m36_10<=m36_10+1;end
else if(m36_10==1250)begin m36_10<=0;io36[10:10]<=~io36[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_11<=149;io36[11:11]<=0;end
else if(m36_11<1250)begin m36_11<=m36_11+1;end
else if(m36_11==1250)begin m36_11<=0;io36[11:11]<=~io36[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_12<=103;io36[12:12]<=0;end
else if(m36_12<1250)begin m36_12<=m36_12+1;end
else if(m36_12==1250)begin m36_12<=0;io36[12:12]<=~io36[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_13<=433;io36[13:13]<=1;end
else if(m36_13<1250)begin m36_13<=m36_13+1;end
else if(m36_13==1250)begin m36_13<=0;io36[13:13]<=~io36[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_14<=274;io36[14:14]<=0;end
else if(m36_14<1250)begin m36_14<=m36_14+1;end
else if(m36_14==1250)begin m36_14<=0;io36[14:14]<=~io36[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_15<=234;io36[15:15]<=0;end
else if(m36_15<1250)begin m36_15<=m36_15+1;end
else if(m36_15==1250)begin m36_15<=0;io36[15:15]<=~io36[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_16<=540;io36[16:16]<=0;end
else if(m36_16<1250)begin m36_16<=m36_16+1;end
else if(m36_16==1250)begin m36_16<=0;io36[16:16]<=~io36[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_17<=90;io36[17:17]<=0;end
else if(m36_17<1250)begin m36_17<=m36_17+1;end
else if(m36_17==1250)begin m36_17<=0;io36[17:17]<=~io36[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_18<=665;io36[18:18]<=1;end
else if(m36_18<1250)begin m36_18<=m36_18+1;end
else if(m36_18==1250)begin m36_18<=0;io36[18:18]<=~io36[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_19<=482;io36[19:19]<=0;end
else if(m36_19<1250)begin m36_19<=m36_19+1;end
else if(m36_19==1250)begin m36_19<=0;io36[19:19]<=~io36[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_20<=148;io36[20:20]<=1;end
else if(m36_20<1250)begin m36_20<=m36_20+1;end
else if(m36_20==1250)begin m36_20<=0;io36[20:20]<=~io36[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_21<=92;io36[21:21]<=1;end
else if(m36_21<1250)begin m36_21<=m36_21+1;end
else if(m36_21==1250)begin m36_21<=0;io36[21:21]<=~io36[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_22<=1221;io36[22:22]<=0;end
else if(m36_22<1250)begin m36_22<=m36_22+1;end
else if(m36_22==1250)begin m36_22<=0;io36[22:22]<=~io36[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_23<=316;io36[23:23]<=0;end
else if(m36_23<1250)begin m36_23<=m36_23+1;end
else if(m36_23==1250)begin m36_23<=0;io36[23:23]<=~io36[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m36_24<=328;io36[24:24]<=1;end
else if(m36_24<1250)begin m36_24<=m36_24+1;end
else if(m36_24==1250)begin m36_24<=0;io36[24:24]<=~io36[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_0<=1052;io37[0:0]<=1;end
else if(m37_0<1250)begin m37_0<=m37_0+1;end
else if(m37_0==1250)begin m37_0<=0;io37[0:0]<=~io37[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_1<=1239;io37[1:1]<=1;end
else if(m37_1<1250)begin m37_1<=m37_1+1;end
else if(m37_1==1250)begin m37_1<=0;io37[1:1]<=~io37[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_2<=927;io37[2:2]<=1;end
else if(m37_2<1250)begin m37_2<=m37_2+1;end
else if(m37_2==1250)begin m37_2<=0;io37[2:2]<=~io37[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_3<=1006;io37[3:3]<=0;end
else if(m37_3<1250)begin m37_3<=m37_3+1;end
else if(m37_3==1250)begin m37_3<=0;io37[3:3]<=~io37[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_4<=849;io37[4:4]<=1;end
else if(m37_4<1250)begin m37_4<=m37_4+1;end
else if(m37_4==1250)begin m37_4<=0;io37[4:4]<=~io37[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_5<=959;io37[5:5]<=0;end
else if(m37_5<1250)begin m37_5<=m37_5+1;end
else if(m37_5==1250)begin m37_5<=0;io37[5:5]<=~io37[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_6<=985;io37[6:6]<=1;end
else if(m37_6<1250)begin m37_6<=m37_6+1;end
else if(m37_6==1250)begin m37_6<=0;io37[6:6]<=~io37[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_7<=624;io37[7:7]<=0;end
else if(m37_7<1250)begin m37_7<=m37_7+1;end
else if(m37_7==1250)begin m37_7<=0;io37[7:7]<=~io37[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_8<=19;io37[8:8]<=1;end
else if(m37_8<1250)begin m37_8<=m37_8+1;end
else if(m37_8==1250)begin m37_8<=0;io37[8:8]<=~io37[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_9<=1138;io37[9:9]<=0;end
else if(m37_9<1250)begin m37_9<=m37_9+1;end
else if(m37_9==1250)begin m37_9<=0;io37[9:9]<=~io37[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_10<=187;io37[10:10]<=0;end
else if(m37_10<1250)begin m37_10<=m37_10+1;end
else if(m37_10==1250)begin m37_10<=0;io37[10:10]<=~io37[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_11<=149;io37[11:11]<=0;end
else if(m37_11<1250)begin m37_11<=m37_11+1;end
else if(m37_11==1250)begin m37_11<=0;io37[11:11]<=~io37[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_12<=103;io37[12:12]<=0;end
else if(m37_12<1250)begin m37_12<=m37_12+1;end
else if(m37_12==1250)begin m37_12<=0;io37[12:12]<=~io37[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_13<=433;io37[13:13]<=1;end
else if(m37_13<1250)begin m37_13<=m37_13+1;end
else if(m37_13==1250)begin m37_13<=0;io37[13:13]<=~io37[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_14<=274;io37[14:14]<=0;end
else if(m37_14<1250)begin m37_14<=m37_14+1;end
else if(m37_14==1250)begin m37_14<=0;io37[14:14]<=~io37[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_15<=234;io37[15:15]<=0;end
else if(m37_15<1250)begin m37_15<=m37_15+1;end
else if(m37_15==1250)begin m37_15<=0;io37[15:15]<=~io37[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_16<=540;io37[16:16]<=0;end
else if(m37_16<1250)begin m37_16<=m37_16+1;end
else if(m37_16==1250)begin m37_16<=0;io37[16:16]<=~io37[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_17<=90;io37[17:17]<=0;end
else if(m37_17<1250)begin m37_17<=m37_17+1;end
else if(m37_17==1250)begin m37_17<=0;io37[17:17]<=~io37[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_18<=665;io37[18:18]<=1;end
else if(m37_18<1250)begin m37_18<=m37_18+1;end
else if(m37_18==1250)begin m37_18<=0;io37[18:18]<=~io37[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_19<=482;io37[19:19]<=0;end
else if(m37_19<1250)begin m37_19<=m37_19+1;end
else if(m37_19==1250)begin m37_19<=0;io37[19:19]<=~io37[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_20<=148;io37[20:20]<=1;end
else if(m37_20<1250)begin m37_20<=m37_20+1;end
else if(m37_20==1250)begin m37_20<=0;io37[20:20]<=~io37[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_21<=92;io37[21:21]<=1;end
else if(m37_21<1250)begin m37_21<=m37_21+1;end
else if(m37_21==1250)begin m37_21<=0;io37[21:21]<=~io37[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_22<=1221;io37[22:22]<=0;end
else if(m37_22<1250)begin m37_22<=m37_22+1;end
else if(m37_22==1250)begin m37_22<=0;io37[22:22]<=~io37[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_23<=316;io37[23:23]<=0;end
else if(m37_23<1250)begin m37_23<=m37_23+1;end
else if(m37_23==1250)begin m37_23<=0;io37[23:23]<=~io37[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m37_24<=328;io37[24:24]<=1;end
else if(m37_24<1250)begin m37_24<=m37_24+1;end
else if(m37_24==1250)begin m37_24<=0;io37[24:24]<=~io37[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_0<=751;io38[0:0]<=0;end
else if(m38_0<1250)begin m38_0<=m38_0+1;end
else if(m38_0==1250)begin m38_0<=0;io38[0:0]<=~io38[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_1<=733;io38[1:1]<=1;end
else if(m38_1<1250)begin m38_1<=m38_1+1;end
else if(m38_1==1250)begin m38_1<=0;io38[1:1]<=~io38[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_2<=721;io38[2:2]<=0;end
else if(m38_2<1250)begin m38_2<=m38_2+1;end
else if(m38_2==1250)begin m38_2<=0;io38[2:2]<=~io38[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_3<=719;io38[3:3]<=1;end
else if(m38_3<1250)begin m38_3<=m38_3+1;end
else if(m38_3==1250)begin m38_3<=0;io38[3:3]<=~io38[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_4<=709;io38[4:4]<=0;end
else if(m38_4<1250)begin m38_4<=m38_4+1;end
else if(m38_4==1250)begin m38_4<=0;io38[4:4]<=~io38[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_5<=825;io38[5:5]<=1;end
else if(m38_5<1250)begin m38_5<=m38_5+1;end
else if(m38_5==1250)begin m38_5<=0;io38[5:5]<=~io38[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_6<=600;io38[6:6]<=0;end
else if(m38_6<1250)begin m38_6<=m38_6+1;end
else if(m38_6==1250)begin m38_6<=0;io38[6:6]<=~io38[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_7<=421;io38[7:7]<=1;end
else if(m38_7<1250)begin m38_7<=m38_7+1;end
else if(m38_7==1250)begin m38_7<=0;io38[7:7]<=~io38[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_8<=607;io38[8:8]<=0;end
else if(m38_8<1250)begin m38_8<=m38_8+1;end
else if(m38_8==1250)begin m38_8<=0;io38[8:8]<=~io38[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_9<=825;io38[9:9]<=1;end
else if(m38_9<1250)begin m38_9<=m38_9+1;end
else if(m38_9==1250)begin m38_9<=0;io38[9:9]<=~io38[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_10<=1227;io38[10:10]<=0;end
else if(m38_10<1250)begin m38_10<=m38_10+1;end
else if(m38_10==1250)begin m38_10<=0;io38[10:10]<=~io38[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_11<=1198;io38[11:11]<=0;end
else if(m38_11<1250)begin m38_11<=m38_11+1;end
else if(m38_11==1250)begin m38_11<=0;io38[11:11]<=~io38[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_12<=1142;io38[12:12]<=0;end
else if(m38_12<1250)begin m38_12<=m38_12+1;end
else if(m38_12==1250)begin m38_12<=0;io38[12:12]<=~io38[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_13<=59;io38[13:13]<=1;end
else if(m38_13<1250)begin m38_13<=m38_13+1;end
else if(m38_13==1250)begin m38_13<=0;io38[13:13]<=~io38[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_14<=5;io38[14:14]<=1;end
else if(m38_14<1250)begin m38_14<=m38_14+1;end
else if(m38_14==1250)begin m38_14<=0;io38[14:14]<=~io38[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_15<=107;io38[15:15]<=1;end
else if(m38_15<1250)begin m38_15<=m38_15+1;end
else if(m38_15==1250)begin m38_15<=0;io38[15:15]<=~io38[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_16<=210;io38[16:16]<=1;end
else if(m38_16<1250)begin m38_16<=m38_16+1;end
else if(m38_16==1250)begin m38_16<=0;io38[16:16]<=~io38[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_17<=1133;io38[17:17]<=0;end
else if(m38_17<1250)begin m38_17<=m38_17+1;end
else if(m38_17==1250)begin m38_17<=0;io38[17:17]<=~io38[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_18<=112;io38[18:18]<=1;end
else if(m38_18<1250)begin m38_18<=m38_18+1;end
else if(m38_18==1250)begin m38_18<=0;io38[18:18]<=~io38[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_19<=169;io38[19:19]<=1;end
else if(m38_19<1250)begin m38_19<=m38_19+1;end
else if(m38_19==1250)begin m38_19<=0;io38[19:19]<=~io38[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_20<=54;io38[20:20]<=0;end
else if(m38_20<1250)begin m38_20<=m38_20+1;end
else if(m38_20==1250)begin m38_20<=0;io38[20:20]<=~io38[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_21<=954;io38[21:21]<=1;end
else if(m38_21<1250)begin m38_21<=m38_21+1;end
else if(m38_21==1250)begin m38_21<=0;io38[21:21]<=~io38[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_22<=1020;io38[22:22]<=1;end
else if(m38_22<1250)begin m38_22<=m38_22+1;end
else if(m38_22==1250)begin m38_22<=0;io38[22:22]<=~io38[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_23<=850;io38[23:23]<=1;end
else if(m38_23<1250)begin m38_23<=m38_23+1;end
else if(m38_23==1250)begin m38_23<=0;io38[23:23]<=~io38[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m38_24<=5;io38[24:24]<=0;end
else if(m38_24<1250)begin m38_24<=m38_24+1;end
else if(m38_24==1250)begin m38_24<=0;io38[24:24]<=~io38[24:24];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_0<=751;io39[0:0]<=0;end
else if(m39_0<1250)begin m39_0<=m39_0+1;end
else if(m39_0==1250)begin m39_0<=0;io39[0:0]<=~io39[0:0];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_1<=733;io39[1:1]<=1;end
else if(m39_1<1250)begin m39_1<=m39_1+1;end
else if(m39_1==1250)begin m39_1<=0;io39[1:1]<=~io39[1:1];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_2<=721;io39[2:2]<=0;end
else if(m39_2<1250)begin m39_2<=m39_2+1;end
else if(m39_2==1250)begin m39_2<=0;io39[2:2]<=~io39[2:2];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_3<=719;io39[3:3]<=1;end
else if(m39_3<1250)begin m39_3<=m39_3+1;end
else if(m39_3==1250)begin m39_3<=0;io39[3:3]<=~io39[3:3];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_4<=709;io39[4:4]<=0;end
else if(m39_4<1250)begin m39_4<=m39_4+1;end
else if(m39_4==1250)begin m39_4<=0;io39[4:4]<=~io39[4:4];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_5<=825;io39[5:5]<=1;end
else if(m39_5<1250)begin m39_5<=m39_5+1;end
else if(m39_5==1250)begin m39_5<=0;io39[5:5]<=~io39[5:5];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_6<=600;io39[6:6]<=0;end
else if(m39_6<1250)begin m39_6<=m39_6+1;end
else if(m39_6==1250)begin m39_6<=0;io39[6:6]<=~io39[6:6];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_7<=421;io39[7:7]<=1;end
else if(m39_7<1250)begin m39_7<=m39_7+1;end
else if(m39_7==1250)begin m39_7<=0;io39[7:7]<=~io39[7:7];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_8<=607;io39[8:8]<=0;end
else if(m39_8<1250)begin m39_8<=m39_8+1;end
else if(m39_8==1250)begin m39_8<=0;io39[8:8]<=~io39[8:8];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_9<=825;io39[9:9]<=1;end
else if(m39_9<1250)begin m39_9<=m39_9+1;end
else if(m39_9==1250)begin m39_9<=0;io39[9:9]<=~io39[9:9];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_10<=1227;io39[10:10]<=0;end
else if(m39_10<1250)begin m39_10<=m39_10+1;end
else if(m39_10==1250)begin m39_10<=0;io39[10:10]<=~io39[10:10];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_11<=1198;io39[11:11]<=0;end
else if(m39_11<1250)begin m39_11<=m39_11+1;end
else if(m39_11==1250)begin m39_11<=0;io39[11:11]<=~io39[11:11];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_12<=1142;io39[12:12]<=0;end
else if(m39_12<1250)begin m39_12<=m39_12+1;end
else if(m39_12==1250)begin m39_12<=0;io39[12:12]<=~io39[12:12];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_13<=59;io39[13:13]<=1;end
else if(m39_13<1250)begin m39_13<=m39_13+1;end
else if(m39_13==1250)begin m39_13<=0;io39[13:13]<=~io39[13:13];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_14<=5;io39[14:14]<=1;end
else if(m39_14<1250)begin m39_14<=m39_14+1;end
else if(m39_14==1250)begin m39_14<=0;io39[14:14]<=~io39[14:14];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_15<=107;io39[15:15]<=1;end
else if(m39_15<1250)begin m39_15<=m39_15+1;end
else if(m39_15==1250)begin m39_15<=0;io39[15:15]<=~io39[15:15];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_16<=210;io39[16:16]<=1;end
else if(m39_16<1250)begin m39_16<=m39_16+1;end
else if(m39_16==1250)begin m39_16<=0;io39[16:16]<=~io39[16:16];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_17<=1133;io39[17:17]<=0;end
else if(m39_17<1250)begin m39_17<=m39_17+1;end
else if(m39_17==1250)begin m39_17<=0;io39[17:17]<=~io39[17:17];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_18<=112;io39[18:18]<=1;end
else if(m39_18<1250)begin m39_18<=m39_18+1;end
else if(m39_18==1250)begin m39_18<=0;io39[18:18]<=~io39[18:18];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_19<=169;io39[19:19]<=1;end
else if(m39_19<1250)begin m39_19<=m39_19+1;end
else if(m39_19==1250)begin m39_19<=0;io39[19:19]<=~io39[19:19];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_20<=54;io39[20:20]<=0;end
else if(m39_20<1250)begin m39_20<=m39_20+1;end
else if(m39_20==1250)begin m39_20<=0;io39[20:20]<=~io39[20:20];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_21<=954;io39[21:21]<=1;end
else if(m39_21<1250)begin m39_21<=m39_21+1;end
else if(m39_21==1250)begin m39_21<=0;io39[21:21]<=~io39[21:21];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_22<=1020;io39[22:22]<=1;end
else if(m39_22<1250)begin m39_22<=m39_22+1;end
else if(m39_22==1250)begin m39_22<=0;io39[22:22]<=~io39[22:22];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_23<=850;io39[23:23]<=1;end
else if(m39_23<1250)begin m39_23<=m39_23+1;end
else if(m39_23==1250)begin m39_23<=0;io39[23:23]<=~io39[23:23];end
end

 always@(posedge clk or posedge reset)
begin
if(reset)begin m39_24<=5;io39[24:24]<=0;end
else if(m39_24<1250)begin m39_24<=m39_24+1;end
else if(m39_24==1250)begin m39_24<=0;io39[24:24]<=~io39[24:24];end
end
